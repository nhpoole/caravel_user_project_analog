magic
tech sky130A
magscale 1 2
timestamp 1624300568
<< pwell >>
rect 294184 -175166 295456 -174946
<< metal1 >>
rect 256482 -91252 256488 -91192
rect 256548 -91252 256760 -91192
rect 274292 -96732 274352 -96726
rect 270862 -96742 270922 -96736
rect 268876 -97882 268882 -97822
rect 268942 -97882 268948 -97822
rect 270862 -98096 270922 -96802
rect 272572 -98078 272578 -98018
rect 272638 -98078 272644 -98018
rect 274292 -98264 274352 -96792
rect 245134 -99510 245140 -99450
rect 245200 -99510 245206 -99450
rect 245140 -101694 245200 -99510
rect 274292 -100226 274352 -100220
rect 269018 -101018 269024 -100958
rect 269084 -101018 269090 -100958
rect 244754 -101754 245200 -101694
rect 274292 -101738 274352 -100286
rect 274294 -103226 274354 -101908
rect 274294 -103292 274354 -103286
rect 272580 -105008 272640 -103626
rect 272580 -105074 272640 -105068
rect 193222 -106070 193370 -106010
rect 193430 -106070 193436 -106010
rect 275244 -107964 275304 -107472
rect 275244 -108030 275304 -108024
rect 243263 -114661 243425 -114603
rect 244188 -114888 244288 -114882
rect 244188 -114994 244288 -114988
rect 340572 -115934 340632 -115928
rect 340632 -115994 341848 -115934
rect 340572 -116000 340632 -115994
rect 206548 -133850 206780 -133844
rect 201482 -134082 206548 -133850
rect 201482 -135136 201542 -134082
rect 206548 -134088 206780 -134082
rect 207072 -133856 207216 -133850
rect 201482 -135196 201624 -135136
rect 199354 -136092 199498 -136086
rect 207072 -136092 207216 -134000
rect 199498 -136236 207216 -136092
rect 207458 -134734 207558 -134728
rect 199354 -136242 199498 -136236
rect 207458 -136628 207558 -134834
rect 207452 -136728 207458 -136628
rect 207558 -136728 207564 -136628
rect 204118 -146250 204124 -146150
rect 204224 -146250 204230 -146150
rect 204124 -148012 204224 -146250
rect 204124 -148118 204224 -148112
rect 195644 -149028 195704 -149022
rect 193666 -149088 195644 -149028
rect 195644 -149094 195704 -149088
rect 259992 -149032 260052 -149026
rect 260052 -149092 260920 -149032
rect 259992 -149098 260052 -149092
rect 340704 -166944 340764 -166938
rect 340764 -167004 341756 -166944
rect 340704 -167010 340764 -167004
rect 339824 -182426 339830 -182366
rect 339890 -182426 339896 -182366
rect 259902 -183556 259962 -183550
rect 184660 -183616 184958 -183556
rect 185018 -183616 185024 -183556
rect 225734 -183616 225954 -183556
rect 226014 -183616 226020 -183556
rect 259962 -183616 260944 -183556
rect 259902 -183622 259962 -183616
rect 339580 -184698 339676 -184692
rect 333766 -184794 333772 -184698
rect 333868 -184794 339580 -184698
rect 339580 -184800 339676 -184794
rect 339678 -184956 339734 -184896
rect 339794 -184956 339800 -184896
rect 334778 -185024 334838 -185018
rect 339830 -185020 339890 -182426
rect 334838 -185084 335058 -185024
rect 339462 -185080 339890 -185020
rect 334778 -185090 334838 -185084
rect 334540 -185242 334636 -185236
rect 334636 -185338 339606 -185242
rect 334540 -185344 334636 -185338
rect 333758 -185882 333764 -185786
rect 333860 -185882 339474 -185786
<< via1 >>
rect 256488 -91252 256548 -91192
rect 270862 -96802 270922 -96742
rect 268882 -97882 268942 -97822
rect 274292 -96792 274352 -96732
rect 272578 -98078 272638 -98018
rect 245140 -99510 245200 -99450
rect 274292 -100286 274352 -100226
rect 269024 -101018 269084 -100958
rect 274294 -103286 274354 -103226
rect 272580 -105068 272640 -105008
rect 193370 -106070 193430 -106010
rect 275244 -108024 275304 -107964
rect 244188 -114988 244288 -114888
rect 340572 -115994 340632 -115934
rect 206548 -134082 206780 -133850
rect 207072 -134000 207216 -133856
rect 199354 -136236 199498 -136092
rect 207458 -134834 207558 -134734
rect 207458 -136728 207558 -136628
rect 204124 -146250 204224 -146150
rect 204124 -148112 204224 -148012
rect 195644 -149088 195704 -149028
rect 259992 -149092 260052 -149032
rect 340704 -167004 340764 -166944
rect 339830 -182426 339890 -182366
rect 184958 -183616 185018 -183556
rect 225954 -183616 226014 -183556
rect 259902 -183616 259962 -183556
rect 333772 -184794 333868 -184698
rect 339580 -184794 339676 -184698
rect 339734 -184956 339794 -184896
rect 334778 -185084 334838 -185024
rect 334540 -185338 334636 -185242
rect 333764 -185882 333860 -185786
<< metal2 >>
rect 199381 -83670 199441 -83504
rect 250374 -91192 256566 -91166
rect 250374 -91252 256488 -91192
rect 256548 -91252 256566 -91192
rect 250374 -91294 256566 -91252
rect 196484 -91585 196584 -91580
rect 196480 -91675 196489 -91585
rect 196579 -91675 196588 -91585
rect 194320 -91947 194420 -91942
rect 194316 -92037 194325 -91947
rect 194415 -92037 194424 -91947
rect 193370 -106010 193430 -106004
rect 193361 -106070 193370 -106010
rect 193430 -106070 193439 -106010
rect 193370 -106076 193430 -106070
rect 194320 -107740 194420 -92037
rect 190376 -107840 194420 -107740
rect 190376 -108711 190476 -107840
rect 190372 -108801 190381 -108711
rect 190471 -108801 190480 -108711
rect 190376 -108806 190476 -108801
rect 196484 -109367 196584 -91675
rect 250374 -92300 250502 -91294
rect 250374 -92437 250502 -92428
rect 266828 -96425 266837 -96291
rect 266971 -96425 266980 -96291
rect 279692 -96386 280120 -96326
rect 265964 -96733 265973 -96567
rect 266139 -96733 266148 -96567
rect 265471 -97957 265480 -97743
rect 265694 -97957 265703 -97743
rect 245104 -99450 262535 -99413
rect 245104 -99510 245140 -99450
rect 245200 -99510 262535 -99450
rect 245104 -99546 262535 -99510
rect 262668 -99546 262677 -99413
rect 265030 -101061 265039 -100911
rect 265189 -101061 265198 -100911
rect 250374 -101205 250502 -101200
rect 250370 -101323 250379 -101205
rect 250497 -101323 250506 -101205
rect 197955 -102432 198015 -102238
rect 198780 -107835 198789 -107705
rect 198919 -107835 198928 -107705
rect 198789 -109177 198919 -107835
rect 210625 -108120 210634 -107984
rect 210770 -108120 210779 -107984
rect 198475 -109307 198919 -109177
rect 196480 -109457 196489 -109367
rect 196579 -109457 196588 -109367
rect 196484 -109462 196584 -109457
rect 191447 -110194 191456 -110134
rect 191516 -110194 191525 -110134
rect 191456 -111380 191516 -110194
rect 194516 -110650 194576 -110641
rect 193494 -110710 194516 -110650
rect 194516 -110719 194576 -110710
rect 191456 -111440 192132 -111380
rect 198475 -112253 198605 -109307
rect 210634 -112248 210770 -108120
rect 211052 -108385 211061 -108259
rect 211187 -108385 211196 -108259
rect 196578 -112346 196790 -112286
rect 196850 -112346 196859 -112286
rect 198471 -112373 198480 -112253
rect 198600 -112373 198609 -112253
rect 208548 -112286 210770 -112248
rect 208476 -112346 210770 -112286
rect 198475 -112378 198605 -112373
rect 208548 -112384 210770 -112346
rect 210170 -114691 210286 -114687
rect 211061 -114691 211187 -108385
rect 211294 -108703 211303 -108569
rect 211437 -108703 211446 -108569
rect 210165 -114696 211187 -114691
rect 210165 -114812 210170 -114696
rect 210286 -114812 211187 -114696
rect 210165 -114817 211187 -114812
rect 210170 -114821 210286 -114817
rect 211303 -115213 211437 -108703
rect 212365 -109046 212374 -108902
rect 212518 -109046 212527 -108902
rect 211557 -114910 211647 -114906
rect 208557 -115250 211437 -115213
rect 196618 -115310 196788 -115250
rect 196848 -115310 196857 -115250
rect 208484 -115310 211437 -115250
rect 208557 -115347 211437 -115310
rect 211552 -114915 211652 -114910
rect 211552 -115005 211557 -114915
rect 211647 -115005 211652 -114915
rect 210524 -115768 210624 -115766
rect 211552 -115768 211652 -115005
rect 210522 -115771 211652 -115768
rect 210520 -115861 210529 -115771
rect 210619 -115861 211652 -115771
rect 210522 -115868 211652 -115861
rect 207458 -120845 207558 -120840
rect 207454 -120935 207463 -120845
rect 207553 -120935 207562 -120845
rect 207063 -121782 207072 -121638
rect 207216 -121782 207225 -121638
rect 206548 -121959 206780 -121954
rect 206544 -122181 206553 -121959
rect 206775 -122181 206784 -121959
rect 206548 -133850 206780 -122181
rect 206542 -134082 206548 -133850
rect 206780 -134082 206786 -133850
rect 207072 -133856 207216 -121782
rect 207066 -134000 207072 -133856
rect 207216 -134000 207222 -133856
rect 207458 -134734 207558 -120935
rect 210524 -122264 210624 -115868
rect 210794 -116871 210894 -116866
rect 210790 -116961 210799 -116871
rect 210889 -116961 210898 -116871
rect 208246 -122364 210624 -122264
rect 207452 -134834 207458 -134734
rect 207558 -134834 207564 -134734
rect 207458 -134838 207558 -134834
rect 195602 -136236 199354 -136092
rect 199498 -136236 199504 -136092
rect 195602 -136441 195746 -136236
rect 195602 -136575 195607 -136441
rect 195741 -136575 195746 -136441
rect 195602 -136580 195746 -136575
rect 195607 -136584 195741 -136580
rect 207458 -136628 207558 -136622
rect 205993 -137496 206083 -137492
rect 207458 -137496 207558 -136728
rect 205988 -137501 207558 -137496
rect 205988 -137591 205993 -137501
rect 206083 -137591 207558 -137501
rect 205988 -137596 207558 -137591
rect 205993 -137600 206083 -137596
rect 204124 -143645 204224 -143640
rect 204120 -143735 204129 -143645
rect 204219 -143735 204228 -143645
rect 204124 -146150 204224 -143735
rect 204811 -144748 204901 -144744
rect 208246 -144748 208346 -122364
rect 204806 -144753 208346 -144748
rect 204806 -144843 204811 -144753
rect 204901 -144843 208346 -144753
rect 204806 -144848 208346 -144843
rect 204811 -144852 204901 -144848
rect 204124 -146256 204224 -146250
rect 158376 -146554 158508 -146518
rect 158376 -146614 160676 -146554
rect 158376 -151698 158508 -146614
rect 204124 -148012 204224 -147992
rect 204118 -148112 204124 -148012
rect 204224 -148112 204230 -148012
rect 195644 -149028 195704 -149019
rect 195638 -149088 195644 -149028
rect 195704 -149088 195710 -149028
rect 195644 -149097 195704 -149088
rect 204124 -153944 204224 -148112
rect 205627 -149274 205717 -149270
rect 210794 -149274 210894 -116961
rect 212374 -121643 212518 -109046
rect 245669 -109410 245678 -109244
rect 245844 -109410 245853 -109244
rect 232501 -109787 232510 -109649
rect 232648 -109787 232657 -109649
rect 218166 -110291 218175 -110141
rect 218325 -110291 218334 -110141
rect 212802 -110527 213034 -110522
rect 212798 -110749 212807 -110527
rect 213029 -110749 213038 -110527
rect 212370 -121777 212379 -121643
rect 212513 -121777 212522 -121643
rect 212374 -121782 212518 -121777
rect 212802 -121954 213034 -110749
rect 212793 -122186 212802 -121954
rect 213034 -122186 213043 -121954
rect 205622 -149279 210896 -149274
rect 205622 -149369 205627 -149279
rect 205717 -149369 210896 -149279
rect 205622 -149374 210896 -149369
rect 205627 -149378 205717 -149374
rect 204124 -154044 210658 -153944
rect 210258 -155363 210267 -155213
rect 210417 -155363 210426 -155213
rect 210036 -169589 210136 -169584
rect 210032 -169679 210041 -169589
rect 210131 -169679 210140 -169589
rect 186411 -183511 186561 -183502
rect 184913 -183556 186411 -183511
rect 184913 -183616 184958 -183556
rect 185018 -183616 186411 -183556
rect 184913 -183661 186411 -183616
rect 186411 -183670 186561 -183661
rect 210036 -184536 210136 -169679
rect 210267 -170068 210417 -155363
rect 210263 -170208 210272 -170068
rect 210412 -170208 210421 -170068
rect 210267 -170213 210417 -170208
rect 210558 -170706 210658 -154044
rect 218175 -155218 218325 -110291
rect 231559 -113926 231568 -113866
rect 231628 -113926 231637 -113866
rect 225357 -114988 225366 -114928
rect 225426 -114988 226682 -114928
rect 225367 -115524 225376 -115464
rect 225436 -115524 226956 -115464
rect 232510 -116116 232648 -109787
rect 244188 -113851 244288 -113846
rect 244184 -113941 244193 -113851
rect 244283 -113941 244292 -113851
rect 244188 -114888 244288 -113941
rect 244182 -114988 244188 -114888
rect 244288 -114988 244294 -114888
rect 231798 -116176 232648 -116116
rect 245678 -116588 245844 -109410
rect 250374 -110560 250502 -101323
rect 264162 -102109 264171 -101963
rect 264317 -102109 264326 -101963
rect 263725 -105406 263734 -105246
rect 263894 -105406 263903 -105246
rect 250365 -110688 250374 -110560
rect 250502 -110688 250511 -110560
rect 250732 -110697 250741 -110539
rect 250899 -110697 250908 -110539
rect 250329 -111474 250338 -111314
rect 250498 -111474 250507 -111314
rect 243378 -116648 245844 -116588
rect 234399 -150312 234522 -150280
rect 234276 -150372 234522 -150312
rect 234399 -151436 234522 -150372
rect 234390 -151559 234399 -151436
rect 234522 -151559 234531 -151436
rect 250338 -151701 250498 -111474
rect 250334 -151851 250343 -151701
rect 250493 -151851 250502 -151701
rect 250338 -151856 250498 -151851
rect 218171 -155358 218180 -155218
rect 218320 -155358 218329 -155218
rect 218175 -155363 218325 -155358
rect 250741 -169266 250899 -110697
rect 255262 -111089 255271 -110943
rect 255417 -111089 255426 -110943
rect 255271 -135621 255417 -111089
rect 263734 -111319 263894 -105406
rect 264171 -110948 264317 -102109
rect 264578 -103529 264587 -103371
rect 264745 -103529 264754 -103371
rect 264587 -110544 264745 -103529
rect 265039 -110146 265189 -101061
rect 265480 -109621 265694 -97957
rect 265973 -109249 266139 -96733
rect 266427 -100176 266436 -100032
rect 266580 -100176 266589 -100032
rect 266436 -108907 266580 -100176
rect 266837 -108574 266971 -96425
rect 274292 -96732 274352 -96723
rect 270862 -96742 270922 -96733
rect 270856 -96802 270862 -96742
rect 270922 -96802 270928 -96742
rect 274286 -96792 274292 -96732
rect 274352 -96792 274358 -96732
rect 274292 -96801 274352 -96792
rect 270862 -96811 270922 -96802
rect 268882 -97822 268942 -97816
rect 268873 -97882 268882 -97822
rect 268942 -97882 268951 -97822
rect 268882 -97888 268942 -97882
rect 272578 -98018 272638 -98009
rect 267503 -98218 267512 -98082
rect 267648 -98218 267657 -98082
rect 272578 -98087 272638 -98078
rect 267190 -98479 267199 -98353
rect 267325 -98479 267334 -98353
rect 267199 -108264 267325 -98479
rect 267512 -107989 267648 -98218
rect 267842 -98312 269144 -98252
rect 267842 -98316 267971 -98312
rect 267841 -107710 267971 -98316
rect 274283 -98418 274294 -98358
rect 274354 -98418 274454 -98358
rect 377155 -99057 377301 -99056
rect 377155 -99117 378347 -99057
rect 268407 -99417 268540 -99411
rect 268403 -99540 268412 -99417
rect 268535 -99540 268544 -99417
rect 268407 -101632 268540 -99540
rect 274292 -100226 274352 -100217
rect 274286 -100286 274292 -100226
rect 274352 -100286 274358 -100226
rect 274292 -100295 274352 -100286
rect 269024 -100958 269084 -100952
rect 269015 -101018 269024 -100958
rect 269084 -101018 269093 -100958
rect 269024 -101024 269084 -101018
rect 268407 -101692 270994 -101632
rect 268136 -101719 268276 -101694
rect 268136 -101809 268161 -101719
rect 268251 -101809 268276 -101719
rect 272569 -101794 272578 -101734
rect 272638 -101794 272816 -101734
rect 268136 -107404 268276 -101809
rect 268882 -101898 269030 -101838
rect 268882 -101998 268942 -101898
rect 268873 -102058 268882 -101998
rect 268942 -102058 268951 -101998
rect 274294 -103226 274354 -103217
rect 274288 -103286 274294 -103226
rect 274354 -103286 274360 -103226
rect 274294 -103295 274354 -103286
rect 279388 -103683 279397 -103533
rect 279547 -103683 279556 -103533
rect 295787 -103572 295796 -103412
rect 295956 -103572 296978 -103412
rect 272580 -105008 272640 -104999
rect 272574 -105068 272580 -105008
rect 272640 -105068 272646 -105008
rect 295832 -105067 296000 -105060
rect 272580 -105077 272640 -105068
rect 275896 -105168 276012 -105108
rect 276072 -105168 276081 -105108
rect 295832 -105205 295849 -105067
rect 295987 -105205 296000 -105067
rect 294183 -107365 294325 -107360
rect 268127 -107544 268136 -107404
rect 268276 -107544 268285 -107404
rect 275792 -107460 276162 -107400
rect 276222 -107460 276231 -107400
rect 294179 -107497 294188 -107365
rect 294320 -107497 294329 -107365
rect 267837 -107830 267846 -107710
rect 267966 -107830 267975 -107710
rect 267841 -107835 267971 -107830
rect 275244 -107964 275304 -107955
rect 267508 -108115 267517 -107989
rect 267643 -108115 267652 -107989
rect 275238 -108024 275244 -107964
rect 275304 -108024 275310 -107964
rect 275244 -108033 275304 -108024
rect 267512 -108120 267648 -108115
rect 275830 -108160 276144 -108100
rect 267195 -108380 267204 -108264
rect 267320 -108380 267329 -108264
rect 267199 -108385 267325 -108380
rect 266833 -108698 266842 -108574
rect 266966 -108698 266975 -108574
rect 266837 -108703 266971 -108698
rect 266432 -109041 266441 -108907
rect 266575 -109041 266584 -108907
rect 266436 -109046 266580 -109041
rect 265969 -109405 265978 -109249
rect 266134 -109405 266143 -109249
rect 265973 -109410 266139 -109405
rect 265476 -109825 265485 -109621
rect 265689 -109825 265698 -109621
rect 265480 -109830 265694 -109825
rect 265035 -110286 265044 -110146
rect 265184 -110286 265193 -110146
rect 265039 -110291 265189 -110286
rect 264583 -110692 264592 -110544
rect 264740 -110692 264749 -110544
rect 264587 -110697 264745 -110692
rect 264167 -111084 264176 -110948
rect 264312 -111084 264321 -110948
rect 264171 -111089 264317 -111084
rect 263730 -111469 263739 -111319
rect 263889 -111469 263898 -111319
rect 263734 -111474 263894 -111469
rect 294183 -124565 294325 -107497
rect 294571 -108186 294717 -108181
rect 294567 -108322 294576 -108186
rect 294712 -108322 294721 -108186
rect 294571 -122067 294717 -108322
rect 294562 -122213 294571 -122067
rect 294717 -122213 294726 -122067
rect 295832 -122978 296000 -105205
rect 296818 -122492 296978 -103572
rect 340522 -115934 340682 -115884
rect 340522 -115994 340572 -115934
rect 340632 -115994 340682 -115934
rect 340080 -118567 340089 -118421
rect 340235 -118567 340244 -118421
rect 297540 -122067 297676 -122063
rect 340089 -122067 340235 -118567
rect 297535 -122072 340235 -122067
rect 297535 -122208 297540 -122072
rect 297676 -122208 340235 -122072
rect 297535 -122213 340235 -122208
rect 297540 -122217 297676 -122213
rect 340522 -122492 340682 -115994
rect 377155 -118426 377301 -99117
rect 384590 -101032 384986 -100972
rect 377792 -101582 378406 -101522
rect 377151 -118562 377160 -118426
rect 377296 -118562 377305 -118426
rect 377155 -118567 377301 -118562
rect 296818 -122652 340682 -122492
rect 295832 -123146 336052 -122978
rect 294183 -124707 295881 -124565
rect 255271 -135767 260089 -135621
rect 259943 -136115 260089 -135767
rect 259943 -136120 260094 -136115
rect 259943 -136256 259953 -136120
rect 260089 -136256 260094 -136120
rect 259943 -136261 260094 -136256
rect 259943 -136265 260089 -136261
rect 294513 -136595 294603 -136586
rect 294513 -136694 294603 -136685
rect 295221 -137023 295230 -136906
rect 295347 -137023 295356 -136906
rect 259992 -149032 260052 -149023
rect 259986 -149092 259992 -149032
rect 260052 -149092 260058 -149032
rect 259992 -149101 260052 -149092
rect 251432 -149386 254490 -149286
rect 258310 -149306 258370 -149297
rect 256528 -149366 258310 -149306
rect 258310 -149375 258370 -149366
rect 250737 -169414 250746 -169266
rect 250894 -169414 250903 -169266
rect 250741 -169419 250899 -169414
rect 210558 -170806 214418 -170706
rect 214318 -179624 214418 -170806
rect 214318 -179684 216972 -179624
rect 227633 -183507 227791 -183498
rect 225905 -183556 227633 -183507
rect 225905 -183616 225954 -183556
rect 226014 -183616 227633 -183556
rect 225905 -183665 227633 -183616
rect 227633 -183674 227791 -183665
rect 251432 -183810 251532 -149386
rect 295230 -150297 295347 -137023
rect 295739 -137257 295881 -124707
rect 298051 -126571 298111 -126488
rect 297116 -126947 297216 -126942
rect 297112 -127037 297121 -126947
rect 297211 -127037 297220 -126947
rect 297116 -136590 297216 -127037
rect 298023 -131005 298140 -126571
rect 297454 -131122 298140 -131005
rect 297107 -136690 297116 -136590
rect 297216 -136690 297225 -136590
rect 297454 -136910 297571 -131122
rect 298051 -135004 298111 -133004
rect 298042 -135064 298051 -135004
rect 298111 -135064 298120 -135004
rect 302051 -135296 302111 -132954
rect 302042 -135356 302051 -135296
rect 302111 -135356 302120 -135296
rect 306051 -135604 306111 -133004
rect 306042 -135664 306051 -135604
rect 306111 -135664 306120 -135604
rect 310051 -135888 310111 -132804
rect 310042 -135948 310051 -135888
rect 310111 -135948 310120 -135888
rect 314051 -136184 314111 -132976
rect 314042 -136244 314051 -136184
rect 314111 -136244 314120 -136184
rect 318051 -136470 318111 -132934
rect 318042 -136530 318051 -136470
rect 318111 -136530 318120 -136470
rect 326051 -136746 326111 -132948
rect 326042 -136806 326051 -136746
rect 326111 -136806 326120 -136746
rect 297453 -137017 297462 -136910
rect 297569 -137017 297578 -136910
rect 297454 -137020 297571 -137017
rect 330051 -137040 330111 -132928
rect 330042 -137100 330051 -137040
rect 330111 -137100 330120 -137040
rect 295739 -137423 334893 -137257
rect 334727 -138572 334893 -137423
rect 334723 -138728 334732 -138572
rect 334888 -138728 334897 -138572
rect 334727 -138733 334893 -138728
rect 253223 -150380 253336 -150377
rect 253218 -150386 253831 -150380
rect 253218 -150499 253223 -150386
rect 253336 -150499 253831 -150386
rect 295221 -150414 295230 -150297
rect 295347 -150414 295356 -150297
rect 253218 -150503 253831 -150499
rect 253223 -150508 253336 -150503
rect 255065 -151856 255074 -151696
rect 255234 -151856 255243 -151696
rect 255074 -170066 255234 -151856
rect 335884 -154082 336052 -123146
rect 336237 -137440 336246 -137340
rect 336346 -137440 336355 -137340
rect 336246 -153801 336346 -137440
rect 377792 -152532 377992 -101582
rect 378162 -137513 378171 -137347
rect 378337 -137513 378346 -137347
rect 378171 -150067 378337 -137513
rect 378171 -150127 378347 -150067
rect 378171 -150180 378337 -150127
rect 384612 -152042 385152 -151982
rect 377792 -152592 378402 -152532
rect 336242 -153891 336251 -153801
rect 336341 -153891 336350 -153801
rect 336246 -153896 336346 -153891
rect 335884 -154250 340818 -154082
rect 340650 -166944 340818 -154250
rect 340650 -167004 340704 -166944
rect 340764 -167004 340818 -166944
rect 340650 -167058 340818 -167004
rect 255074 -170226 260016 -170066
rect 259856 -170776 260016 -170226
rect 377792 -170574 377992 -152592
rect 259854 -170808 260016 -170776
rect 260014 -170968 260016 -170808
rect 259854 -170974 260016 -170968
rect 340100 -170656 340210 -170644
rect 340100 -170716 340116 -170656
rect 340176 -170716 340210 -170656
rect 259854 -170977 260014 -170974
rect 294346 -175096 294530 -175036
rect 294590 -175096 294599 -175036
rect 299029 -178252 299038 -178192
rect 299098 -178252 299192 -178192
rect 334540 -180252 334636 -180243
rect 259902 -183556 259962 -183547
rect 259896 -183616 259902 -183556
rect 259962 -183616 259968 -183556
rect 259902 -183625 259962 -183616
rect 251432 -183830 254488 -183810
rect 258292 -183830 258352 -183821
rect 251432 -183890 254562 -183830
rect 256782 -183890 258292 -183830
rect 251432 -183910 254488 -183890
rect 258292 -183899 258352 -183890
rect 210027 -184636 210036 -184536
rect 210136 -184636 210145 -184536
rect 173363 -184718 173506 -184705
rect 173138 -184778 173506 -184718
rect 173363 -186046 173506 -184778
rect 253275 -184880 253284 -184760
rect 253404 -184880 253413 -184760
rect 253284 -184938 253404 -184880
rect 253284 -184998 253882 -184938
rect 253284 -185028 253404 -184998
rect 173359 -186179 173368 -186046
rect 173501 -186179 173510 -186046
rect 173363 -186183 173506 -186179
rect 298051 -186346 298111 -184146
rect 298042 -186406 298051 -186346
rect 298111 -186406 298120 -186346
rect 302051 -186638 302111 -184096
rect 302042 -186698 302051 -186638
rect 302111 -186698 302120 -186638
rect 306051 -186946 306111 -184146
rect 306042 -187006 306051 -186946
rect 306111 -187006 306120 -186946
rect 310051 -187230 310111 -183946
rect 310042 -187290 310051 -187230
rect 310111 -187290 310120 -187230
rect 314051 -187526 314111 -184118
rect 314042 -187586 314051 -187526
rect 314111 -187586 314120 -187526
rect 318051 -187812 318111 -184076
rect 318042 -187872 318051 -187812
rect 318111 -187872 318120 -187812
rect 326051 -188088 326111 -184090
rect 326042 -188148 326051 -188088
rect 326111 -188148 326120 -188088
rect 330051 -188382 330111 -184070
rect 333772 -184698 333868 -184692
rect 333763 -184794 333772 -184698
rect 333868 -184794 333877 -184698
rect 333772 -184800 333868 -184794
rect 334540 -185242 334636 -180348
rect 339830 -182366 339890 -182360
rect 338791 -182426 338800 -182366
rect 338860 -182426 339830 -182366
rect 339830 -182432 339890 -182426
rect 339574 -184794 339580 -184698
rect 339676 -184794 339682 -184698
rect 334737 -185024 334880 -184982
rect 334737 -185084 334778 -185024
rect 334838 -185084 334880 -185024
rect 334534 -185338 334540 -185242
rect 334636 -185338 334642 -185242
rect 333764 -185786 333860 -185780
rect 333755 -185882 333764 -185786
rect 333860 -185882 333869 -185786
rect 333764 -185888 333860 -185882
rect 334737 -186042 334880 -185084
rect 339580 -185466 339676 -184794
rect 339734 -184896 339794 -184890
rect 340100 -184896 340210 -170716
rect 377783 -170774 377792 -170574
rect 377992 -170774 378001 -170574
rect 339794 -184956 340210 -184896
rect 339734 -184962 339794 -184956
rect 334728 -186185 334737 -186042
rect 334880 -186185 334889 -186042
rect 330042 -188442 330051 -188382
rect 330111 -188442 330120 -188382
<< via2 >>
rect 196489 -91675 196579 -91585
rect 194325 -92037 194415 -91947
rect 193370 -106070 193430 -106010
rect 190381 -108801 190471 -108711
rect 250374 -92428 250502 -92300
rect 266837 -96425 266971 -96291
rect 265973 -96733 266139 -96567
rect 265480 -97957 265694 -97743
rect 262535 -99546 262668 -99413
rect 265039 -101061 265189 -100911
rect 250379 -101323 250497 -101205
rect 198789 -107835 198919 -107705
rect 210634 -108120 210770 -107984
rect 196489 -109457 196579 -109367
rect 191456 -110194 191516 -110134
rect 194516 -110710 194576 -110650
rect 211061 -108385 211187 -108259
rect 196790 -112346 196850 -112286
rect 198480 -112373 198600 -112253
rect 211303 -108703 211437 -108569
rect 210170 -114812 210286 -114696
rect 212374 -109046 212518 -108902
rect 196788 -115310 196848 -115250
rect 211557 -115005 211647 -114915
rect 210529 -115861 210619 -115771
rect 207463 -120935 207553 -120845
rect 207072 -121782 207216 -121638
rect 206553 -122181 206775 -121959
rect 210799 -116961 210889 -116871
rect 195607 -136575 195741 -136441
rect 205993 -137591 206083 -137501
rect 204129 -143735 204219 -143645
rect 204811 -144843 204901 -144753
rect 195644 -149088 195704 -149028
rect 245678 -109410 245844 -109244
rect 232510 -109787 232648 -109649
rect 218175 -110291 218325 -110141
rect 212807 -110749 213029 -110527
rect 212379 -121777 212513 -121643
rect 212802 -122186 213034 -121954
rect 205627 -149369 205717 -149279
rect 210267 -155363 210417 -155213
rect 210041 -169679 210131 -169589
rect 186411 -183661 186561 -183511
rect 210272 -170208 210412 -170068
rect 231568 -113926 231628 -113866
rect 225366 -114988 225426 -114928
rect 225376 -115524 225436 -115464
rect 244193 -113941 244283 -113851
rect 264171 -102109 264317 -101963
rect 263734 -105406 263894 -105246
rect 250374 -110688 250502 -110560
rect 250741 -110697 250899 -110539
rect 250338 -111474 250498 -111314
rect 234399 -151559 234522 -151436
rect 250343 -151851 250493 -151701
rect 218180 -155358 218320 -155218
rect 255271 -111089 255417 -110943
rect 264587 -103529 264745 -103371
rect 266436 -100176 266580 -100032
rect 270862 -96802 270922 -96742
rect 274292 -96792 274352 -96732
rect 268882 -97882 268942 -97822
rect 272578 -98078 272638 -98018
rect 267512 -98218 267648 -98082
rect 267199 -98479 267325 -98353
rect 274294 -98418 274354 -98358
rect 268412 -99540 268535 -99417
rect 274292 -100286 274352 -100226
rect 269024 -101018 269084 -100958
rect 268161 -101809 268251 -101719
rect 272578 -101794 272638 -101734
rect 268882 -102058 268942 -101998
rect 274294 -103286 274354 -103226
rect 279397 -103683 279547 -103533
rect 295796 -103572 295956 -103412
rect 272580 -105068 272640 -105008
rect 276012 -105168 276072 -105108
rect 295849 -105205 295987 -105067
rect 268136 -107544 268276 -107404
rect 276162 -107460 276222 -107400
rect 294188 -107497 294320 -107365
rect 267846 -107830 267966 -107710
rect 267517 -108115 267643 -107989
rect 275244 -108024 275304 -107964
rect 267204 -108380 267320 -108264
rect 266842 -108698 266966 -108574
rect 266441 -109041 266575 -108907
rect 265978 -109405 266134 -109249
rect 265485 -109825 265689 -109621
rect 265044 -110286 265184 -110146
rect 264592 -110692 264740 -110544
rect 264176 -111084 264312 -110948
rect 263739 -111469 263889 -111319
rect 294576 -108322 294712 -108186
rect 294571 -122213 294717 -122067
rect 340089 -118567 340235 -118421
rect 297540 -122208 297676 -122072
rect 377160 -118562 377296 -118426
rect 259953 -136256 260089 -136120
rect 294513 -136685 294603 -136595
rect 295230 -137023 295347 -136906
rect 259992 -149092 260052 -149032
rect 258310 -149366 258370 -149306
rect 250746 -169414 250894 -169266
rect 227633 -183665 227791 -183507
rect 297121 -127037 297211 -126947
rect 297116 -136690 297216 -136590
rect 298051 -135064 298111 -135004
rect 302051 -135356 302111 -135296
rect 306051 -135664 306111 -135604
rect 310051 -135948 310111 -135888
rect 314051 -136244 314111 -136184
rect 318051 -136530 318111 -136470
rect 326051 -136806 326111 -136746
rect 297462 -137017 297569 -136910
rect 330051 -137100 330111 -137040
rect 334732 -138728 334888 -138572
rect 253223 -150499 253336 -150386
rect 295230 -150414 295347 -150297
rect 255074 -151856 255234 -151696
rect 336246 -137440 336346 -137340
rect 378171 -137513 378337 -137347
rect 336251 -153891 336341 -153801
rect 259854 -170968 260014 -170808
rect 340116 -170716 340176 -170656
rect 294530 -175096 294590 -175036
rect 299038 -178252 299098 -178192
rect 334540 -180348 334636 -180252
rect 259902 -183616 259962 -183556
rect 258292 -183890 258352 -183830
rect 210036 -184636 210136 -184536
rect 253284 -184880 253404 -184760
rect 173368 -186179 173501 -186046
rect 298051 -186406 298111 -186346
rect 302051 -186698 302111 -186638
rect 306051 -187006 306111 -186946
rect 310051 -187290 310111 -187230
rect 314051 -187586 314111 -187526
rect 318051 -187872 318111 -187812
rect 326051 -188148 326111 -188088
rect 333772 -184794 333868 -184698
rect 338800 -182426 338860 -182366
rect 333764 -185882 333860 -185786
rect 377792 -170774 377992 -170574
rect 334737 -186185 334880 -186042
rect 330051 -188442 330111 -188382
<< metal3 >>
rect 196370 -91585 196584 -91580
rect 196370 -91675 196489 -91585
rect 196579 -91675 196584 -91585
rect 196370 -91680 196584 -91675
rect 194320 -91947 194420 -91942
rect 194320 -92037 194325 -91947
rect 194415 -92037 194420 -91947
rect 194320 -92042 194420 -92037
rect 250369 -92300 250507 -92295
rect 250369 -92428 250374 -92300
rect 250502 -92428 250507 -92300
rect 250369 -92433 250507 -92428
rect 200736 -99558 201006 -99458
rect 250374 -101205 250502 -92433
rect 266832 -96291 266976 -96286
rect 266832 -96425 266837 -96291
rect 266971 -96295 266976 -96291
rect 266971 -96425 274386 -96295
rect 266832 -96430 266976 -96425
rect 265968 -96567 266144 -96562
rect 265968 -96733 265973 -96567
rect 266139 -96580 266144 -96567
rect 266139 -96726 270968 -96580
rect 266139 -96733 266144 -96726
rect 265968 -96738 266144 -96733
rect 270822 -96742 270968 -96726
rect 270822 -96802 270862 -96742
rect 270922 -96802 270968 -96742
rect 270822 -96826 270968 -96802
rect 274256 -96732 274386 -96425
rect 274256 -96792 274292 -96732
rect 274352 -96792 274386 -96732
rect 274256 -96816 274386 -96792
rect 265475 -97743 265699 -97738
rect 265475 -97957 265480 -97743
rect 265694 -97782 265699 -97743
rect 265694 -97822 268974 -97782
rect 265694 -97882 268882 -97822
rect 268942 -97882 268974 -97822
rect 265694 -97922 268974 -97882
rect 265694 -97957 265699 -97922
rect 265475 -97962 265699 -97957
rect 272541 -98018 272671 -97995
rect 267507 -98082 267653 -98077
rect 267507 -98218 267512 -98082
rect 267648 -98086 267653 -98082
rect 272541 -98078 272578 -98018
rect 272638 -98078 272671 -98018
rect 272541 -98086 272671 -98078
rect 267648 -98216 272671 -98086
rect 267648 -98218 267653 -98216
rect 267507 -98223 267653 -98218
rect 267194 -98352 267330 -98348
rect 267194 -98353 274356 -98352
rect 267194 -98479 267199 -98353
rect 267325 -98358 274359 -98353
rect 267325 -98418 274294 -98358
rect 274354 -98418 274359 -98358
rect 267325 -98423 274359 -98418
rect 267325 -98476 274356 -98423
rect 267325 -98479 267330 -98476
rect 267194 -98484 267330 -98479
rect 262530 -99412 262673 -99408
rect 262530 -99413 268540 -99412
rect 262530 -99546 262535 -99413
rect 262668 -99417 268540 -99413
rect 262668 -99540 268412 -99417
rect 268535 -99540 268540 -99417
rect 262668 -99545 268540 -99540
rect 262668 -99546 262673 -99545
rect 262530 -99551 262673 -99546
rect 266431 -100030 266585 -100027
rect 266431 -100032 274378 -100030
rect 266431 -100176 266436 -100032
rect 266580 -100144 274378 -100032
rect 266580 -100176 266585 -100144
rect 266431 -100181 266585 -100176
rect 274264 -100226 274378 -100144
rect 274264 -100286 274292 -100226
rect 274352 -100286 274378 -100226
rect 274264 -100298 274378 -100286
rect 257354 -100828 257834 -100728
rect 265034 -100911 265194 -100906
rect 265034 -101061 265039 -100911
rect 265189 -100914 265194 -100911
rect 265189 -100958 269112 -100914
rect 265189 -101018 269024 -100958
rect 269084 -101018 269112 -100958
rect 265189 -101061 269112 -101018
rect 265034 -101064 269112 -101061
rect 265034 -101066 265194 -101064
rect 250374 -101323 250379 -101205
rect 250497 -101323 250502 -101205
rect 250374 -101328 250502 -101323
rect 268156 -101719 272660 -101714
rect 268156 -101809 268161 -101719
rect 268251 -101734 272660 -101719
rect 268251 -101794 272578 -101734
rect 272638 -101794 272660 -101734
rect 268251 -101809 272660 -101794
rect 268156 -101814 272660 -101809
rect 264166 -101962 264322 -101958
rect 264166 -101963 268970 -101962
rect 264166 -102109 264171 -101963
rect 264317 -101998 268970 -101963
rect 264317 -102058 268882 -101998
rect 268942 -102058 268970 -101998
rect 264317 -102109 268970 -102058
rect 264166 -102110 268970 -102109
rect 264166 -102114 264322 -102110
rect 274254 -103226 274400 -103192
rect 274254 -103286 274294 -103226
rect 274354 -103286 274400 -103226
rect 264582 -103371 264750 -103366
rect 264582 -103529 264587 -103371
rect 264745 -103375 264750 -103371
rect 274254 -103375 274400 -103286
rect 264745 -103521 274400 -103375
rect 295791 -103412 295961 -103407
rect 264745 -103529 264750 -103521
rect 264582 -103534 264750 -103529
rect 279392 -103533 295796 -103412
rect 279392 -103683 279397 -103533
rect 279547 -103572 295796 -103533
rect 295956 -103572 295961 -103412
rect 279547 -103683 279552 -103572
rect 295791 -103577 295961 -103572
rect 279392 -103688 279552 -103683
rect 272530 -105008 272686 -104986
rect 272530 -105068 272580 -105008
rect 272640 -105068 272686 -105008
rect 263729 -105246 263899 -105241
rect 257776 -105356 258178 -105256
rect 263729 -105406 263734 -105246
rect 263894 -105250 263899 -105246
rect 272530 -105250 272686 -105068
rect 275988 -105067 295992 -105062
rect 275988 -105108 295849 -105067
rect 275988 -105168 276012 -105108
rect 276072 -105168 295849 -105108
rect 275988 -105205 295849 -105168
rect 295987 -105205 295992 -105067
rect 275988 -105210 295992 -105205
rect 263894 -105406 272686 -105250
rect 263729 -105411 263899 -105406
rect 193330 -106010 197124 -105970
rect 193330 -106070 193370 -106010
rect 193430 -106070 197124 -106010
rect 193330 -106110 197124 -106070
rect 196984 -107404 197124 -106110
rect 276138 -107365 294325 -107360
rect 268131 -107404 268281 -107399
rect 196984 -107544 268136 -107404
rect 268276 -107544 268281 -107404
rect 276138 -107400 294188 -107365
rect 276138 -107460 276162 -107400
rect 276222 -107460 294188 -107400
rect 276138 -107497 294188 -107460
rect 294320 -107497 294325 -107365
rect 276138 -107502 294325 -107497
rect 268131 -107549 268281 -107544
rect 198784 -107705 198924 -107700
rect 198784 -107835 198789 -107705
rect 198919 -107710 267971 -107705
rect 198919 -107830 267846 -107710
rect 267966 -107830 267971 -107710
rect 198919 -107835 267971 -107830
rect 198784 -107840 198924 -107835
rect 275204 -107964 275350 -107944
rect 210629 -107984 210775 -107979
rect 210629 -108120 210634 -107984
rect 210770 -107989 267648 -107984
rect 210770 -108115 267517 -107989
rect 267643 -108115 267648 -107989
rect 210770 -108120 267648 -108115
rect 275204 -108024 275244 -107964
rect 275304 -108024 275350 -107964
rect 210629 -108125 210775 -108120
rect 275204 -108181 275350 -108024
rect 275204 -108186 294717 -108181
rect 211056 -108259 211192 -108254
rect 211056 -108385 211061 -108259
rect 211187 -108264 267325 -108259
rect 211187 -108380 267204 -108264
rect 267320 -108380 267325 -108264
rect 275204 -108322 294576 -108186
rect 294712 -108322 294717 -108186
rect 275204 -108327 294717 -108322
rect 211187 -108385 267325 -108380
rect 211056 -108390 211192 -108385
rect 211298 -108569 211442 -108564
rect 211298 -108703 211303 -108569
rect 211437 -108574 266971 -108569
rect 211437 -108698 266842 -108574
rect 266966 -108698 266971 -108574
rect 211437 -108703 266971 -108698
rect 190376 -108711 190476 -108706
rect 211298 -108708 211442 -108703
rect 190376 -108801 190381 -108711
rect 190471 -108801 190476 -108711
rect 190376 -110116 190476 -108801
rect 212369 -108902 212523 -108897
rect 212369 -109046 212374 -108902
rect 212518 -108907 266580 -108902
rect 212518 -109041 266441 -108907
rect 266575 -109041 266580 -108907
rect 212518 -109046 266580 -109041
rect 212369 -109051 212523 -109046
rect 245673 -109244 245849 -109239
rect 196484 -109367 196584 -109362
rect 196484 -109457 196489 -109367
rect 196579 -109457 196584 -109367
rect 245673 -109410 245678 -109244
rect 245844 -109249 266139 -109244
rect 245844 -109405 265978 -109249
rect 266134 -109405 266139 -109249
rect 245844 -109410 266139 -109405
rect 245673 -109415 245849 -109410
rect 196484 -110116 196584 -109457
rect 232508 -109621 265694 -109616
rect 232508 -109644 265485 -109621
rect 232505 -109649 265485 -109644
rect 232505 -109787 232510 -109649
rect 232648 -109787 265485 -109649
rect 232505 -109792 265485 -109787
rect 232508 -109825 265485 -109792
rect 265689 -109825 265694 -109621
rect 232508 -109830 265694 -109825
rect 190376 -110134 191542 -110116
rect 190376 -110194 191456 -110134
rect 191516 -110194 191542 -110134
rect 190376 -110216 191542 -110194
rect 194496 -110216 196584 -110116
rect 218170 -110141 218330 -110136
rect 194496 -110650 194596 -110216
rect 218170 -110291 218175 -110141
rect 218325 -110146 265189 -110141
rect 218325 -110286 265044 -110146
rect 265184 -110286 265189 -110146
rect 218325 -110291 265189 -110286
rect 218170 -110296 218330 -110291
rect 194496 -110710 194516 -110650
rect 194576 -110710 194596 -110650
rect 194496 -110732 194596 -110710
rect 212802 -110527 250536 -110522
rect 212802 -110749 212807 -110527
rect 213029 -110560 250536 -110527
rect 213029 -110688 250374 -110560
rect 250502 -110688 250536 -110560
rect 213029 -110749 250536 -110688
rect 250736 -110539 250904 -110534
rect 250736 -110697 250741 -110539
rect 250899 -110544 264745 -110539
rect 250899 -110692 264592 -110544
rect 264740 -110692 264745 -110544
rect 250899 -110697 264745 -110692
rect 250736 -110702 250904 -110697
rect 212802 -110754 250536 -110749
rect 255266 -110943 255422 -110938
rect 255266 -111089 255271 -110943
rect 255417 -110948 264317 -110943
rect 255417 -111084 264176 -110948
rect 264312 -111084 264317 -110948
rect 255417 -111089 264317 -111084
rect 255266 -111094 255422 -111089
rect 336284 -111122 336606 -111022
rect 250333 -111314 250503 -111309
rect 250333 -111474 250338 -111314
rect 250498 -111319 263894 -111314
rect 250498 -111469 263739 -111319
rect 263889 -111469 263894 -111319
rect 250498 -111474 263894 -111469
rect 250333 -111479 250503 -111474
rect 186620 -111908 186720 -111614
rect 186882 -111772 186982 -111506
rect 196756 -112253 198605 -112248
rect 196756 -112286 198480 -112253
rect 196756 -112346 196790 -112286
rect 196850 -112346 198480 -112286
rect 196756 -112373 198480 -112346
rect 198600 -112373 198605 -112253
rect 196756 -112378 198605 -112373
rect 231546 -113851 244288 -113846
rect 231546 -113866 244193 -113851
rect 231546 -113926 231568 -113866
rect 231628 -113926 244193 -113866
rect 231546 -113941 244193 -113926
rect 244283 -113941 244288 -113851
rect 231546 -113946 244288 -113941
rect 199111 -114696 210291 -114691
rect 199111 -114812 210170 -114696
rect 210286 -114812 210291 -114696
rect 199111 -114817 210291 -114812
rect 199111 -115218 199237 -114817
rect 211552 -114915 225442 -114910
rect 211552 -115005 211557 -114915
rect 211647 -114928 225442 -114915
rect 211647 -114988 225366 -114928
rect 225426 -114988 225442 -114928
rect 211647 -115005 225442 -114988
rect 211552 -115010 225442 -115005
rect 196754 -115250 199237 -115218
rect 196754 -115310 196788 -115250
rect 196848 -115310 199237 -115250
rect 196754 -115344 199237 -115310
rect 210808 -115464 225456 -115442
rect 210808 -115524 225376 -115464
rect 225436 -115524 225456 -115464
rect 210808 -115542 225456 -115524
rect 210524 -115771 210624 -115644
rect 210524 -115861 210529 -115771
rect 210619 -115861 210624 -115771
rect 210524 -115866 210624 -115861
rect 206496 -117378 206596 -116016
rect 210794 -116871 210894 -116692
rect 210794 -116961 210799 -116871
rect 210889 -116961 210894 -116871
rect 210794 -116966 210894 -116961
rect 206496 -117478 207558 -117378
rect 207458 -120845 207558 -117478
rect 340084 -118421 340240 -118416
rect 340084 -118567 340089 -118421
rect 340235 -118426 377301 -118421
rect 340235 -118562 377160 -118426
rect 377296 -118562 377301 -118426
rect 340235 -118567 377301 -118562
rect 340084 -118572 340240 -118567
rect 338785 -119638 338885 -119002
rect 207458 -120935 207463 -120845
rect 207553 -120935 207558 -120845
rect 207458 -120940 207558 -120935
rect 207067 -121638 207221 -121633
rect 207067 -121782 207072 -121638
rect 207216 -121643 212518 -121638
rect 207216 -121777 212379 -121643
rect 212513 -121777 212518 -121643
rect 207216 -121782 212518 -121777
rect 207067 -121787 207221 -121782
rect 212797 -121954 213039 -121949
rect 206548 -121959 212802 -121954
rect 206548 -122181 206553 -121959
rect 206775 -122181 212802 -121959
rect 206548 -122186 212802 -122181
rect 213034 -122186 213039 -121954
rect 212797 -122191 213039 -122186
rect 294566 -122067 294722 -122062
rect 294566 -122213 294571 -122067
rect 294717 -122072 297681 -122067
rect 294717 -122208 297540 -122072
rect 297676 -122208 297681 -122072
rect 294717 -122213 297681 -122208
rect 294566 -122218 294722 -122213
rect 338785 -124480 338885 -123906
rect 338785 -124586 338885 -124580
rect 297116 -126947 298230 -126942
rect 297116 -127037 297121 -126947
rect 297211 -127037 298230 -126947
rect 297116 -127042 298230 -127037
rect 297550 -132004 297938 -131904
rect 297746 -133988 298290 -133888
rect 298030 -135004 336458 -134982
rect 298030 -135064 298051 -135004
rect 298111 -135064 336458 -135004
rect 298030 -135082 336458 -135064
rect 302028 -135296 336456 -135274
rect 302028 -135356 302051 -135296
rect 302111 -135356 336456 -135296
rect 302028 -135374 336456 -135356
rect 306032 -135604 336464 -135584
rect 306032 -135664 306051 -135604
rect 306111 -135664 336464 -135604
rect 306032 -135684 336464 -135664
rect 310030 -135888 336472 -135868
rect 310030 -135948 310051 -135888
rect 310111 -135948 336472 -135888
rect 310030 -135968 336472 -135948
rect 259948 -136120 260094 -136115
rect 259948 -136256 259953 -136120
rect 260089 -136256 260094 -136120
rect 195602 -136441 195746 -136436
rect 195602 -136575 195607 -136441
rect 195741 -136575 195746 -136441
rect 195602 -149028 195746 -136575
rect 203960 -137501 206088 -137496
rect 203960 -137591 205993 -137501
rect 206083 -137591 206088 -137501
rect 203960 -137596 206088 -137591
rect 204124 -143641 204224 -143640
rect 204119 -143739 204125 -143641
rect 204223 -143739 204229 -143641
rect 204124 -143740 204224 -143739
rect 204348 -144753 204906 -144748
rect 204348 -144843 204811 -144753
rect 204901 -144843 204906 -144753
rect 204348 -144848 204906 -144843
rect 195602 -149088 195644 -149028
rect 195704 -149088 195746 -149028
rect 195602 -149116 195746 -149088
rect 259948 -149032 260094 -136256
rect 314026 -136184 336470 -136166
rect 314026 -136244 314051 -136184
rect 314111 -136244 336470 -136184
rect 314026 -136266 336470 -136244
rect 318028 -136470 336472 -136448
rect 318028 -136530 318051 -136470
rect 318111 -136530 336472 -136470
rect 318028 -136548 336472 -136530
rect 297111 -136590 297221 -136585
rect 294508 -136595 297116 -136590
rect 294508 -136685 294513 -136595
rect 294603 -136685 297116 -136595
rect 294508 -136690 297116 -136685
rect 297216 -136690 297221 -136590
rect 297111 -136695 297221 -136690
rect 326026 -136746 336488 -136726
rect 326026 -136806 326051 -136746
rect 326111 -136806 336488 -136746
rect 326026 -136826 336488 -136806
rect 295225 -136905 295352 -136901
rect 295225 -136906 297574 -136905
rect 295225 -137023 295230 -136906
rect 295347 -136910 297574 -136906
rect 295347 -137017 297462 -136910
rect 297569 -137017 297574 -136910
rect 295347 -137022 297574 -137017
rect 295347 -137023 295352 -137022
rect 295225 -137028 295352 -137023
rect 330026 -137040 336500 -137020
rect 330026 -137100 330051 -137040
rect 330111 -137100 336500 -137040
rect 330026 -137120 336500 -137100
rect 336241 -137340 336351 -137335
rect 336241 -137440 336246 -137340
rect 336346 -137342 336351 -137340
rect 338786 -137342 338884 -137337
rect 336346 -137343 338885 -137342
rect 336346 -137440 338786 -137343
rect 336241 -137441 338786 -137440
rect 338884 -137441 338885 -137343
rect 378166 -137347 378342 -137342
rect 336241 -137442 338885 -137441
rect 336241 -137445 336351 -137442
rect 338786 -137447 338884 -137442
rect 351353 -137513 378171 -137347
rect 378337 -137513 378342 -137347
rect 351353 -138567 351519 -137513
rect 378166 -137518 378342 -137513
rect 334727 -138572 351519 -138567
rect 334727 -138728 334732 -138572
rect 334888 -138728 351519 -138572
rect 334727 -138733 351519 -138728
rect 259948 -149092 259992 -149032
rect 260052 -149092 260094 -149032
rect 259948 -149118 260094 -149092
rect 203784 -149279 205722 -149274
rect 203784 -149369 205627 -149279
rect 205717 -149369 205722 -149279
rect 203784 -149374 205722 -149369
rect 258292 -149306 258409 -149262
rect 258292 -149366 258310 -149306
rect 258370 -149366 258409 -149306
rect 258292 -150296 258409 -149366
rect 295225 -150296 295352 -150292
rect 258292 -150297 295352 -150296
rect 253218 -150386 253341 -150381
rect 253218 -150499 253223 -150386
rect 253336 -150499 253341 -150386
rect 258292 -150413 295230 -150297
rect 295225 -150414 295230 -150413
rect 295347 -150414 295352 -150297
rect 295225 -150419 295352 -150414
rect 234394 -151435 234527 -151431
rect 253218 -151435 253341 -150499
rect 234394 -151436 253341 -151435
rect 234394 -151559 234399 -151436
rect 234522 -151558 253341 -151436
rect 234522 -151559 234527 -151558
rect 234394 -151564 234527 -151559
rect 255069 -151696 255239 -151691
rect 250338 -151701 255074 -151696
rect 250338 -151851 250343 -151701
rect 250493 -151851 255074 -151701
rect 250338 -151856 255074 -151851
rect 255234 -151856 255239 -151696
rect 255069 -151861 255239 -151856
rect 336246 -153801 336346 -153796
rect 336246 -153891 336251 -153801
rect 336341 -153891 336346 -153801
rect 210262 -155213 210422 -155208
rect 210262 -155363 210267 -155213
rect 210417 -155218 218325 -155213
rect 210417 -155358 218180 -155218
rect 218320 -155358 218325 -155218
rect 210417 -155363 218325 -155358
rect 210262 -155368 210422 -155363
rect 336246 -161489 336346 -153891
rect 336241 -161587 336247 -161489
rect 336345 -161587 336351 -161489
rect 336246 -161588 336346 -161587
rect 336364 -162132 336720 -162032
rect 338785 -166628 338885 -166622
rect 338785 -167752 338885 -166728
rect 227633 -169266 250899 -169261
rect 227633 -169414 250746 -169266
rect 250894 -169414 250899 -169266
rect 227633 -169419 250899 -169414
rect 187545 -169584 187643 -169579
rect 187544 -169585 210136 -169584
rect 187544 -169683 187545 -169585
rect 187643 -169589 210136 -169585
rect 187643 -169679 210041 -169589
rect 210131 -169679 210136 -169589
rect 187643 -169683 210136 -169679
rect 187544 -169684 210136 -169683
rect 187545 -169689 187643 -169684
rect 186411 -170068 210417 -170063
rect 186411 -170208 210272 -170068
rect 210412 -170208 210417 -170068
rect 186411 -170213 210417 -170208
rect 186411 -183506 186561 -170213
rect 227633 -183502 227791 -169419
rect 377787 -170574 377997 -170569
rect 340092 -170656 377792 -170574
rect 340092 -170716 340116 -170656
rect 340176 -170716 377792 -170656
rect 340092 -170774 377792 -170716
rect 377992 -170774 377997 -170574
rect 377787 -170779 377997 -170774
rect 259849 -170808 260019 -170803
rect 259849 -170968 259854 -170808
rect 260014 -170968 260019 -170808
rect 259849 -170973 260019 -170968
rect 186406 -183511 186566 -183506
rect 186406 -183661 186411 -183511
rect 186561 -183661 186566 -183511
rect 186406 -183666 186566 -183661
rect 227628 -183507 227796 -183502
rect 227628 -183665 227633 -183507
rect 227791 -183665 227796 -183507
rect 259854 -183556 260014 -170973
rect 294506 -175036 295272 -175012
rect 294506 -175096 294530 -175036
rect 294590 -175096 295272 -175036
rect 294506 -175112 295272 -175096
rect 295172 -177952 295272 -175112
rect 295172 -178052 298374 -177952
rect 259854 -183616 259902 -183556
rect 259962 -183616 260014 -183556
rect 259854 -183646 260014 -183616
rect 296002 -178192 299114 -178170
rect 296002 -178252 299038 -178192
rect 299098 -178252 299114 -178192
rect 296002 -178270 299114 -178252
rect 227628 -183670 227796 -183665
rect 258272 -183830 258372 -183802
rect 258272 -183890 258292 -183830
rect 258352 -183890 258372 -183830
rect 210031 -184536 210141 -184531
rect 210031 -184636 210036 -184536
rect 210136 -184636 211630 -184536
rect 210031 -184641 210141 -184636
rect 211530 -184760 211630 -184636
rect 253279 -184760 253409 -184755
rect 211530 -184880 253284 -184760
rect 253404 -184880 253409 -184760
rect 253279 -184885 253409 -184880
rect 258272 -184818 258372 -183890
rect 296002 -184818 296102 -178270
rect 334535 -180247 334641 -180241
rect 334535 -180348 334540 -180343
rect 334636 -180348 334641 -180343
rect 334535 -180353 334641 -180348
rect 338785 -182366 338885 -175208
rect 338785 -182426 338800 -182366
rect 338860 -182426 338885 -182366
rect 338785 -182438 338885 -182426
rect 297634 -183014 298016 -182914
rect 333761 -184799 333767 -184693
rect 333863 -184698 333873 -184693
rect 333868 -184794 333873 -184698
rect 333863 -184799 333873 -184794
rect 258272 -184918 296102 -184818
rect 297882 -184998 298348 -184898
rect 333753 -185887 333759 -185781
rect 333855 -185786 333865 -185781
rect 333860 -185882 333865 -185786
rect 333855 -185887 333865 -185882
rect 334732 -186041 334885 -186037
rect 173363 -186042 334885 -186041
rect 173363 -186046 334737 -186042
rect 173363 -186179 173368 -186046
rect 173501 -186179 334737 -186046
rect 173363 -186184 334737 -186179
rect 334732 -186185 334737 -186184
rect 334880 -186185 334885 -186042
rect 334732 -186190 334885 -186185
rect 298030 -186346 336458 -186324
rect 298030 -186406 298051 -186346
rect 298111 -186406 336458 -186346
rect 298030 -186424 336458 -186406
rect 302028 -186638 336456 -186616
rect 302028 -186698 302051 -186638
rect 302111 -186698 336456 -186638
rect 302028 -186716 336456 -186698
rect 306032 -186946 336464 -186926
rect 306032 -187006 306051 -186946
rect 306111 -187006 336464 -186946
rect 306032 -187026 336464 -187006
rect 310030 -187230 336472 -187210
rect 310030 -187290 310051 -187230
rect 310111 -187290 336472 -187230
rect 310030 -187310 336472 -187290
rect 314026 -187526 336470 -187508
rect 314026 -187586 314051 -187526
rect 314111 -187586 336470 -187526
rect 314026 -187608 336470 -187586
rect 318028 -187812 336472 -187790
rect 318028 -187872 318051 -187812
rect 318111 -187872 336472 -187812
rect 318028 -187890 336472 -187872
rect 326026 -188088 336488 -188068
rect 326026 -188148 326051 -188088
rect 326111 -188148 336488 -188088
rect 326026 -188168 336488 -188148
rect 330026 -188382 336500 -188362
rect 330026 -188442 330051 -188382
rect 330111 -188442 336500 -188382
rect 330026 -188462 336500 -188442
<< via3 >>
rect 338785 -124580 338885 -124480
rect 204125 -143645 204223 -143641
rect 204125 -143735 204129 -143645
rect 204129 -143735 204219 -143645
rect 204219 -143735 204223 -143645
rect 204125 -143739 204223 -143735
rect 338786 -137441 338884 -137343
rect 336247 -161587 336345 -161489
rect 338785 -166728 338885 -166628
rect 187545 -169683 187643 -169585
rect 334535 -180252 334641 -180247
rect 334535 -180343 334540 -180252
rect 334540 -180343 334636 -180252
rect 334636 -180343 334641 -180252
rect 333767 -184698 333863 -184693
rect 333767 -184794 333772 -184698
rect 333772 -184794 333863 -184698
rect 333767 -184799 333863 -184794
rect 333759 -185786 333855 -185781
rect 333759 -185882 333764 -185786
rect 333764 -185882 333855 -185786
rect 333759 -185887 333855 -185882
<< metal4 >>
rect 157844 -78376 160852 -78352
rect 157844 -79128 157868 -78376
rect 158620 -79128 160852 -78376
rect 157844 -79152 160852 -79128
rect 247146 -79140 295982 -78340
rect 280914 -96106 295976 -95306
rect 258602 -107340 269368 -106540
rect 158644 -108980 187308 -108180
rect 268534 -109174 269368 -107340
rect 268534 -109208 269334 -109174
rect 229772 -112180 236238 -111508
rect 208338 -113420 212086 -113396
rect 208338 -114172 211310 -113420
rect 212062 -114172 212086 -113420
rect 208338 -114196 212086 -114172
rect 225610 -118458 236324 -117514
rect 342116 -118218 384856 -117418
rect 190842 -118958 208773 -118846
rect 185684 -119740 208773 -118958
rect 185684 -120184 185708 -119740
rect 186460 -120184 208773 -119740
rect 190842 -120512 208773 -120184
rect 247830 -119074 250970 -118274
rect 250052 -120516 256954 -119716
rect 293920 -120516 295980 -119716
rect 210357 -125412 222055 -123602
rect 296768 -124076 302270 -123388
rect 338784 -124480 338886 -124479
rect 338784 -124580 338785 -124480
rect 338885 -124580 338886 -124480
rect 338784 -124581 338886 -124580
rect 295296 -129556 302212 -128756
rect 296776 -134888 301586 -134200
rect 338785 -137343 338885 -124581
rect 338785 -137441 338786 -137343
rect 338884 -137441 338885 -137343
rect 338785 -137442 338885 -137441
rect 204124 -143641 204224 -141788
rect 210437 -143414 221791 -141512
rect 204124 -143739 204125 -143641
rect 204223 -143739 204224 -143641
rect 204124 -143740 204224 -143739
rect 200065 -151312 221000 -150512
rect 247926 -150538 261544 -150516
rect 247926 -151290 250952 -150538
rect 251704 -151290 261544 -150538
rect 247926 -151316 261544 -151290
rect 380500 -154034 384852 -153234
rect 249184 -154278 256746 -154240
rect 249184 -155030 249300 -154278
rect 250052 -155030 256746 -154278
rect 249184 -155040 256746 -155030
rect 293878 -155040 295976 -154240
rect 336246 -161489 338885 -161488
rect 336246 -161587 336247 -161489
rect 336345 -161587 338885 -161489
rect 336246 -161588 338885 -161587
rect 338785 -166627 338885 -161588
rect 338784 -166628 338886 -166627
rect 338784 -166728 338785 -166628
rect 338885 -166728 338886 -166628
rect 338784 -166729 338886 -166728
rect 186884 -169585 187644 -169584
rect 186884 -169683 187545 -169585
rect 187643 -169683 187644 -169585
rect 186884 -169684 187644 -169683
rect 296776 -175086 301464 -174398
rect 297398 -180566 302070 -179766
rect 334534 -180247 334642 -180246
rect 334534 -180343 334535 -180247
rect 334641 -180343 334642 -180247
rect 334534 -180344 334642 -180343
rect 333766 -184693 333864 -184692
rect 333766 -184799 333767 -184693
rect 333863 -184799 333864 -184693
rect 333766 -184800 333864 -184799
rect 247432 -185840 250928 -185040
rect 251728 -185840 258624 -185040
rect 295308 -185060 297398 -185036
rect 295308 -185812 296622 -185060
rect 297374 -185812 297398 -185060
rect 295308 -185836 297398 -185812
rect 333758 -185781 333856 -185780
rect 333758 -185887 333759 -185781
rect 333855 -185887 333856 -185781
rect 333758 -185888 333856 -185887
<< via4 >>
rect 157868 -79128 158620 -78376
rect 295982 -79140 296782 -78340
rect 295976 -96106 296776 -95306
rect 211286 -107340 212086 -106540
rect 250952 -107316 251704 -106564
rect 157844 -108980 158644 -108180
rect 211310 -114172 212062 -113420
rect 384856 -118218 385656 -117418
rect 185708 -120492 186460 -119740
rect 208773 -120512 210439 -118846
rect 250970 -119074 251770 -118274
rect 249252 -120516 250052 -119716
rect 295980 -120516 296780 -119716
rect 208547 -125412 210357 -123602
rect 296080 -124076 296768 -123388
rect 294496 -129556 295296 -128756
rect 296088 -134888 296776 -134200
rect 208535 -143414 210437 -141512
rect 250952 -151290 251704 -150538
rect 294520 -151322 295272 -150570
rect 384852 -154034 385652 -153234
rect 249300 -155030 250052 -154278
rect 295976 -155040 296776 -154240
rect 296088 -175086 296776 -174398
rect 296598 -180566 297398 -179766
rect 250928 -185840 251728 -185040
rect 296622 -185812 297374 -185060
<< metal5 >>
rect 296088 -78316 296776 -78314
rect 295958 -78340 296806 -78316
rect 157844 -78376 158644 -78352
rect 157844 -79128 157868 -78376
rect 158620 -79128 158644 -78376
rect 157844 -108156 158644 -79128
rect 295958 -79140 295982 -78340
rect 296782 -79140 296806 -78340
rect 295958 -79164 296806 -79140
rect 296088 -95282 296776 -79164
rect 295952 -95306 296800 -95282
rect 295952 -96106 295976 -95306
rect 296776 -96106 296800 -95306
rect 295952 -96130 296800 -96106
rect 211262 -106540 212110 -106516
rect 211262 -107340 211286 -106540
rect 212086 -107340 212110 -106540
rect 211262 -107364 212110 -107340
rect 250928 -106564 251728 -106540
rect 250928 -107316 250952 -106564
rect 251704 -107316 251728 -106564
rect 157820 -108180 158668 -108156
rect 157820 -108980 157844 -108180
rect 158644 -108980 158668 -108180
rect 157820 -109004 158668 -108980
rect 211286 -113420 212086 -107364
rect 211286 -114172 211310 -113420
rect 212062 -114172 212086 -113420
rect 211286 -114196 212086 -114172
rect 185684 -119740 186484 -117842
rect 250928 -118250 251728 -107316
rect 250928 -118274 251794 -118250
rect 185684 -120492 185708 -119740
rect 186460 -120492 186484 -119740
rect 185684 -120516 186484 -120492
rect 208535 -118822 210437 -118641
rect 208535 -118846 210463 -118822
rect 208535 -120512 208773 -118846
rect 210439 -120512 210463 -118846
rect 250928 -119074 250970 -118274
rect 251770 -119074 251794 -118274
rect 250928 -119098 251794 -119074
rect 208535 -120536 210463 -120512
rect 249228 -119716 250076 -119692
rect 249228 -120516 249252 -119716
rect 250052 -120516 250076 -119716
rect 208535 -123578 210437 -120536
rect 249228 -120540 250076 -120516
rect 208523 -123602 210437 -123578
rect 208523 -125412 208547 -123602
rect 210357 -125412 210437 -123602
rect 208523 -125436 210437 -125412
rect 208535 -141488 210437 -125436
rect 250928 -135242 251728 -119098
rect 296088 -119692 296776 -96130
rect 384832 -117418 385680 -117394
rect 384832 -118218 384856 -117418
rect 385656 -118218 385680 -117418
rect 384832 -118242 385680 -118218
rect 295956 -119716 296804 -119692
rect 295956 -120516 295980 -119716
rect 296780 -120516 296804 -119716
rect 295956 -120540 296804 -120516
rect 296088 -123364 296776 -120540
rect 296056 -123388 296792 -123364
rect 296056 -124076 296080 -123388
rect 296768 -124076 296792 -123388
rect 296056 -124100 296792 -124076
rect 294472 -128756 295320 -128732
rect 294472 -129556 294496 -128756
rect 295296 -129556 295320 -128756
rect 294472 -129580 295320 -129556
rect 250928 -136042 256670 -135242
rect 208511 -141512 210461 -141488
rect 208511 -143414 208535 -141512
rect 210437 -143414 210461 -141512
rect 208511 -143438 210461 -143414
rect 249276 -154278 250076 -149618
rect 249276 -155030 249300 -154278
rect 250052 -155030 250076 -154278
rect 249276 -155054 250076 -155030
rect 250928 -150538 251728 -136042
rect 250928 -151290 250952 -150538
rect 251704 -151290 251728 -150538
rect 250928 -185016 251728 -151290
rect 294496 -150570 295296 -129580
rect 296088 -134176 296776 -124100
rect 296064 -134200 296800 -134176
rect 296064 -134888 296088 -134200
rect 296776 -134888 296800 -134200
rect 296064 -134912 296800 -134888
rect 294496 -151322 294520 -150570
rect 295272 -151322 295296 -150570
rect 294496 -151346 295296 -151322
rect 296088 -154216 296776 -134912
rect 335069 -139430 335869 -122300
rect 384852 -153210 385652 -118242
rect 384828 -153234 385676 -153210
rect 384828 -154034 384852 -153234
rect 385652 -154034 385676 -153234
rect 384828 -154058 385676 -154034
rect 295952 -154240 296800 -154216
rect 295952 -155040 295976 -154240
rect 296776 -155040 296800 -154240
rect 295952 -155064 296800 -155040
rect 296088 -174374 296776 -155064
rect 296064 -174398 296800 -174374
rect 296064 -175086 296088 -174398
rect 296776 -175086 296800 -174398
rect 296064 -175110 296800 -175086
rect 296574 -179766 297422 -179742
rect 296574 -180566 296598 -179766
rect 297398 -180566 297422 -179766
rect 296574 -180590 297422 -180566
rect 250904 -185040 251752 -185016
rect 250904 -185840 250928 -185040
rect 251728 -185840 251752 -185040
rect 296598 -185060 297398 -180590
rect 296598 -185812 296622 -185060
rect 297374 -185812 297398 -185060
rect 296598 -185836 297398 -185812
rect 250904 -185864 251752 -185840
use peak_detector  peak_detector_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/peak_detector
timestamp 1624298412
transform 1 0 173892 0 1 -185010
box -16568 -888 76950 30794
use biquad_gm_c_filter  biquad_gm_c_filter_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/biquad_gm_c_filter
timestamp 1624298412
transform 1 0 187212 0 1 -113396
box -1552 -6022 23682 5240
use sample_and_hold  sample_and_hold_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/sample_and_hold
timestamp 1624298412
transform 1 0 253730 0 1 -149196
box -1766 -2178 42040 29480
use sample_and_hold  sample_and_hold_1
timestamp 1624298412
transform 1 0 253730 0 1 -183720
box -1766 -2178 42040 29480
use comparator  comparator_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/continuous_time_comparator
timestamp 1624298412
transform 1 0 229012 0 1 -114708
box -3400 -3600 3400 3200
use diff_to_se_converter  diff_to_se_converter_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_to_se_converter
timestamp 1624300568
transform -1 0 194530 0 1 -150652
box -13514 -718 35912 30940
use input_amplifier  input_amplifier_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/input_amplifier
timestamp 1624300568
transform -1 0 248960 0 1 -106680
box -13477 -718 90192 28340
use low_freq_pll  low_freq_pll_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/low_freq_pll
timestamp 1624300568
transform 1 0 211340 0 1 -129086
box 7294 -22262 38743 17578
use bias_current_distribution  bias_current_distribution_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/bias_current_distribution
timestamp 1624298412
transform 1 0 268974 0 1 -98308
box -440 -10900 12700 3000
use dac_8bit  dac_8bit_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/dac_8bit
timestamp 1624300568
transform 1 0 326281 0 1 -59040
box -29235 -75848 58525 12
use dac_8bit  dac_8bit_1
timestamp 1624300568
transform 1 0 326281 0 1 -110050
box -29235 -75848 58525 12
use pulse_generator  pulse_generator_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/pulse_generator
timestamp 1624300568
transform -1 0 339666 0 1 -185362
box -72 -526 4688 670
<< labels >>
flabel via4 251350 -185504 251356 -185498 1 FreeSans 480 0 0 0 VSS
flabel metal4 252560 -154626 252626 -154538 1 FreeSans 480 0 0 0 VDD
flabel metal3 336386 -135042 336406 -135028 1 FreeSans 480 0 0 0 q7A
flabel metal3 336392 -135326 336404 -135314 1 FreeSans 480 0 0 0 q6A
flabel metal3 336398 -135642 336402 -135632 1 FreeSans 480 0 0 0 q5A
flabel metal3 336394 -135924 336410 -135904 1 FreeSans 480 0 0 0 q4A
flabel metal3 336392 -136230 336400 -136218 1 FreeSans 480 0 0 0 q3A
flabel metal3 336402 -136498 336418 -136486 1 FreeSans 480 0 0 0 q2A
flabel metal3 336410 -136792 336422 -136778 1 FreeSans 480 0 0 0 q1A
flabel metal3 336388 -137080 336412 -137056 1 FreeSans 480 0 0 0 q0A
flabel metal3 297672 -182972 297684 -182956 1 FreeSans 480 0 0 0 vlowB
flabel metal3 297928 -184958 297938 -184946 1 FreeSans 480 0 0 0 vrefB
flabel metal3 297592 -131956 297600 -131944 1 FreeSans 480 0 0 0 vlowA
flabel metal3 297816 -133942 297832 -133926 1 FreeSans 480 0 0 0 vrefA
flabel metal2 377876 -131602 377900 -131586 1 FreeSans 480 0 0 0 adc_clk
flabel metal3 336360 -186390 336394 -186356 1 FreeSans 480 0 0 0 q7B
flabel metal3 336352 -186674 336380 -186650 1 FreeSans 480 0 0 0 q6B
flabel metal3 336360 -187004 336384 -186976 1 FreeSans 480 0 0 0 q5B
flabel metal3 336346 -187278 336366 -187250 1 FreeSans 480 0 0 0 q4B
flabel metal3 336360 -187572 336380 -187544 1 FreeSans 480 0 0 0 q3B
flabel metal3 336360 -187860 336384 -187828 1 FreeSans 480 0 0 0 q2B
flabel metal3 336380 -188130 336404 -188102 1 FreeSans 480 0 0 0 q1B
flabel metal3 336376 -188428 336404 -188404 1 FreeSans 480 0 0 0 q0B
flabel metal2 340136 -184296 340154 -184284 1 FreeSans 480 0 0 0 adc_clk
flabel metal1 339852 -184050 339870 -184034 1 FreeSans 480 0 0 0 sample
flabel metal3 296034 -178004 296042 -178000 1 FreeSans 480 0 0 0 vpeak_sampled
flabel metal2 297150 -127600 297164 -127580 1 FreeSans 480 0 0 0 vcp_sampled
flabel metal3 252684 -184830 252706 -184802 1 FreeSans 480 0 0 0 vpeak
flabel metal3 252302 -151498 252314 -151468 1 FreeSans 480 0 0 0 vcp
flabel metal3 233848 -113906 233872 -113882 1 FreeSans 480 0 0 0 vcomp
flabel metal2 207498 -136864 207514 -136850 1 FreeSans 480 0 0 0 vocm_filt
flabel metal2 190664 -107802 190678 -107782 1 FreeSans 480 0 0 0 vampp
flabel metal2 210568 -116246 210592 -116228 1 FreeSans 480 0 0 0 vfiltp
flabel metal2 210828 -117166 210854 -117146 1 FreeSans 480 0 0 0 vfiltm
flabel metal3 186922 -111650 186936 -111624 1 FreeSans 480 0 0 0 vintm
flabel metal3 186656 -111776 186678 -111748 1 FreeSans 480 0 0 0 vintp
flabel metal2 197976 -102334 197986 -102326 1 FreeSans 480 0 0 0 gain_ctrl_0
flabel metal3 200836 -99526 200866 -99496 1 FreeSans 480 0 0 0 vocm
flabel metal2 204160 -152696 204176 -152670 1 FreeSans 480 0 0 0 vse
flabel metal2 276048 -108136 276068 -108126 1 FreeSans 480 0 0 0 vbiasn
flabel metal2 280014 -96358 280028 -96342 1 FreeSans 480 0 0 0 vbiasp
flabel metal3 336424 -111070 336442 -111054 1 FreeSans 480 0 0 0 adc_vcaparrayA
flabel metal3 336538 -162098 336560 -162076 1 FreeSans 480 0 0 0 adc_vcaparrayB
flabel metal2 384914 -101012 384932 -101002 1 FreeSans 480 0 0 0 adc_compA
flabel metal2 384800 -152028 384810 -152024 1 FreeSans 480 0 0 0 adc_compB
flabel metal2 196520 -107834 196534 -107828 1 FreeSans 480 0 0 0 vampm
flabel metal2 199398 -83588 199416 -83576 1 FreeSans 480 0 0 0 gain_ctrl_1
flabel metal2 334794 -185540 334800 -185524 1 FreeSans 480 0 0 0 peak_detector_rst
flabel metal2 256268 -91234 256286 -91216 1 FreeSans 480 0 0 0 rst_n
flabel metal3 257576 -100770 257584 -100760 1 FreeSans 480 0 0 0 vhpf
flabel metal3 257954 -105312 257972 -105298 1 FreeSans 480 0 0 0 vincm
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nwell >>
rect 74185 58186 76094 59026
<< pwell >>
rect 76043 58128 76073 58130
rect 76043 57472 76094 58128
<< viali >>
rect 74267 58956 74487 58990
rect 75759 58956 75961 58990
rect 74219 58320 74257 58892
rect 75995 58318 76031 58894
rect 74267 58222 74487 58256
rect 75759 58224 75961 58258
rect 76164 58116 76212 58164
rect 76268 58146 76314 58186
rect 74291 58020 74499 58058
rect 75763 58022 75961 58060
rect 74219 57604 74255 57960
rect 75995 57604 76033 57960
rect 74289 57508 74497 57544
rect 75761 57506 75963 57542
<< metal1 >>
rect 74208 59056 76044 59116
rect 74208 59004 74268 59056
rect 74319 59004 74379 59056
rect 74208 59002 74379 59004
rect 74453 59002 74513 59056
rect 74208 58990 74513 59002
rect 74208 58956 74267 58990
rect 74487 58956 74513 58990
rect 74208 58942 74513 58956
rect 74208 58892 74269 58942
rect 74208 58862 74219 58892
rect 74209 58634 74219 58862
rect 74208 58574 74219 58634
rect 74209 58320 74219 58574
rect 74257 58634 74269 58892
rect 74319 58634 74379 58942
rect 74453 58851 74513 58942
rect 74709 59008 74769 59009
rect 75485 59008 75545 59014
rect 74709 58948 75485 59008
rect 74709 58853 74769 58948
rect 74967 58851 75027 58948
rect 75225 58853 75285 58948
rect 75485 58853 75545 58948
rect 75741 59006 75801 59056
rect 75869 59006 75929 59056
rect 75984 59006 76044 59056
rect 75741 58990 76044 59006
rect 75741 58956 75759 58990
rect 75961 58956 76044 58990
rect 75741 58942 76044 58956
rect 75741 58851 75801 58942
rect 74257 58574 74379 58634
rect 75869 58636 75929 58942
rect 75983 58894 76044 58942
rect 75983 58636 75995 58894
rect 75869 58576 75995 58636
rect 74257 58320 74269 58574
rect 74209 58270 74269 58320
rect 74321 58270 74381 58452
rect 74449 58270 74509 58358
rect 74208 58256 74509 58270
rect 74208 58222 74267 58256
rect 74487 58222 74509 58256
rect 74208 58210 74509 58222
rect 74579 58093 74639 58463
rect 74837 58242 74897 58438
rect 74831 58182 74837 58242
rect 74897 58182 74903 58242
rect 74207 58058 74511 58068
rect 74207 58020 74291 58058
rect 74499 58020 74511 58058
rect 74573 58033 74579 58093
rect 74639 58033 74645 58093
rect 74207 58008 74511 58020
rect 74207 57960 74267 58008
rect 74207 57604 74219 57960
rect 74255 57604 74267 57960
rect 74321 57820 74381 58008
rect 74451 57920 74511 58008
rect 74579 57833 74639 58033
rect 74837 57900 74897 58182
rect 75095 58093 75155 58461
rect 75355 58242 75415 58456
rect 75349 58182 75355 58242
rect 75415 58182 75421 58242
rect 75089 58033 75095 58093
rect 75155 58033 75161 58093
rect 74837 57834 74899 57900
rect 74207 57555 74267 57604
rect 74323 57555 74383 57733
rect 74839 57654 74899 57834
rect 75095 57714 75155 58033
rect 75355 57654 75415 58182
rect 75613 58093 75673 58461
rect 75737 58270 75797 58358
rect 75871 58270 75931 58448
rect 75983 58318 75995 58576
rect 76031 58878 76044 58894
rect 76031 58518 76043 58878
rect 76031 58422 76144 58518
rect 76031 58318 76043 58422
rect 75983 58270 76043 58318
rect 75737 58258 76043 58270
rect 75737 58224 75759 58258
rect 75961 58224 76043 58258
rect 75737 58210 76043 58224
rect 76476 58192 76536 58198
rect 76256 58186 76476 58192
rect 76158 58170 76218 58176
rect 76152 58110 76158 58170
rect 76218 58110 76224 58170
rect 76256 58146 76268 58186
rect 76314 58146 76476 58186
rect 76256 58132 76476 58146
rect 76476 58126 76536 58132
rect 76158 58104 76218 58110
rect 75613 57831 75673 58033
rect 75743 58060 76045 58070
rect 75743 58022 75763 58060
rect 75961 58022 76045 58060
rect 75743 58010 76045 58022
rect 75743 57922 75803 58010
rect 75871 57824 75931 58010
rect 75985 57974 76045 58010
rect 75985 57960 76136 57974
rect 74451 57555 74511 57644
rect 74207 57544 74511 57555
rect 74207 57508 74289 57544
rect 74497 57508 74511 57544
rect 74207 57495 74511 57508
rect 74207 57438 74267 57495
rect 74208 57420 74267 57438
rect 74323 57420 74383 57495
rect 74451 57420 74511 57495
rect 74709 57545 74769 57645
rect 74969 57545 75029 57645
rect 75227 57545 75287 57643
rect 75483 57545 75543 57643
rect 75741 57555 75801 57646
rect 75869 57555 75929 57727
rect 75985 57604 75995 57960
rect 76033 57878 76136 57960
rect 76033 57604 76045 57878
rect 75985 57555 76045 57604
rect 74709 57485 75483 57545
rect 75543 57485 75549 57545
rect 75741 57542 76045 57555
rect 75741 57506 75761 57542
rect 75963 57506 76045 57542
rect 75741 57495 76045 57506
rect 75741 57420 75801 57495
rect 75869 57420 75929 57495
rect 75985 57420 76045 57495
rect 74208 57360 76046 57420
<< via1 >>
rect 75485 58948 75545 59008
rect 74837 58182 74897 58242
rect 74579 58033 74639 58093
rect 75355 58182 75415 58242
rect 75095 58033 75155 58093
rect 76158 58164 76218 58170
rect 76158 58116 76164 58164
rect 76164 58116 76212 58164
rect 76212 58116 76218 58164
rect 76158 58110 76218 58116
rect 76476 58132 76536 58192
rect 75613 58033 75673 58093
rect 75483 57485 75543 57545
<< metal2 >>
rect 75479 58948 75485 59008
rect 75545 58948 76144 59008
rect 74837 58242 74897 58248
rect 75355 58242 75415 58248
rect 74897 58182 75355 58242
rect 74837 58176 74897 58182
rect 75355 58176 75415 58182
rect 76084 58170 76144 58948
rect 76084 58110 76158 58170
rect 76218 58110 76224 58170
rect 76470 58132 76476 58192
rect 76536 58132 76542 58192
rect 74579 58093 74639 58099
rect 75095 58093 75155 58099
rect 74568 58033 74579 58093
rect 74639 58033 75095 58093
rect 75155 58033 75613 58093
rect 75673 58033 75679 58093
rect 74579 58027 74639 58033
rect 75095 58027 75155 58033
rect 75483 57545 75543 57551
rect 76476 57546 76536 58132
rect 75990 57545 76536 57546
rect 75543 57486 76536 57545
rect 75543 57485 76094 57486
rect 75483 57479 75543 57485
use sky130_fd_pr__nfet_01v8_N6QVV6  sky130_fd_pr__nfet_01v8_N6QVV6_0
timestamp 1623971255
transform 1 0 75126 0 1 57782
box -941 -310 941 310
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623971255
transform -1 0 76381 0 1 57926
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_hvt_SCHXZ7  sky130_fd_pr__pfet_01v8_hvt_SCHXZ7_0
timestamp 1623971255
transform 1 0 75126 0 1 58606
box -941 -419 941 419
<< labels >>
flabel metal1 76416 58154 76424 58160 1 FreeSans 480 0 0 0 tx
flabel metal1 74598 58134 74608 58142 1 FreeSans 480 0 0 0 out
flabel metal1 74860 58140 74870 58148 1 FreeSans 480 0 0 0 in
flabel metal1 75114 59082 75124 59092 1 FreeSans 480 0 0 0 VDD
flabel metal1 75112 57392 75120 57398 1 FreeSans 480 0 0 0 VSS
flabel metal2 76114 58656 76124 58664 1 FreeSans 480 0 0 0 txb
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nmos >>
rect -100 -200 100 200
<< ndiff >>
rect -158 188 -100 200
rect -158 -188 -146 188
rect -112 -188 -100 188
rect -158 -200 -100 -188
rect 100 188 158 200
rect 100 -188 112 188
rect 146 -188 158 188
rect 100 -200 158 -188
<< ndiffc >>
rect -146 -188 -112 188
rect 112 -188 146 188
<< poly >>
rect -66 272 66 288
rect -66 255 -50 272
rect -100 238 -50 255
rect 50 255 66 272
rect 50 238 100 255
rect -100 200 100 238
rect -100 -238 100 -200
rect -100 -255 -50 -238
rect -66 -272 -50 -255
rect 50 -255 100 -238
rect 50 -272 66 -255
rect -66 -288 66 -272
<< polycont >>
rect -50 238 50 272
rect -50 -272 50 -238
<< locali >>
rect -66 238 -50 272
rect 50 238 66 272
rect -146 188 -112 204
rect -146 -204 -112 -188
rect 112 188 146 204
rect 112 -204 146 -188
rect -66 -272 -50 -238
rect 50 -272 66 -238
<< viali >>
rect -42 238 42 272
rect -146 -188 -112 188
rect 112 -188 146 188
rect -42 -272 42 -238
<< metal1 >>
rect -54 272 54 278
rect -54 238 -42 272
rect 42 238 54 272
rect -54 232 54 238
rect -152 188 -106 200
rect -152 -188 -146 188
rect -112 -188 -106 188
rect -152 -200 -106 -188
rect 106 188 152 200
rect 106 -188 112 188
rect 146 -188 152 188
rect 106 -200 152 -188
rect -54 -238 54 -232
rect -54 -272 -42 -238
rect 42 -272 54 -238
rect -54 -278 54 -272
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 2 l 1 m 1 nf 1 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>

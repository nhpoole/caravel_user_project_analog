magic
tech sky130A
magscale 1 2
timestamp 1623984492
<< nwell >>
rect -2562 -664 6962 2702
<< pwell >>
rect -2558 -3818 6960 -720
<< psubdiff >>
rect -2522 -1618 -2360 -1518
rect 6760 -1618 6922 -1518
rect -2522 -1680 -2422 -1618
rect -2522 -3682 -2422 -3620
rect 6822 -1680 6922 -1618
rect 6822 -3682 6922 -3620
rect -2522 -3782 -2360 -3682
rect 6760 -3782 6922 -3682
<< nsubdiff >>
rect -2522 2562 -2360 2662
rect 6760 2562 6922 2662
rect -2522 2500 -2422 2562
rect -2522 458 -2422 520
rect 6822 2500 6922 2562
rect 6822 458 6922 520
rect -2522 358 -2360 458
rect 6760 358 6922 458
<< psubdiffcont >>
rect -2360 -1618 6760 -1518
rect -2522 -3620 -2422 -1680
rect 6822 -3620 6922 -1680
rect -2360 -3782 6760 -3682
<< nsubdiffcont >>
rect -2360 2562 6760 2662
rect -2522 520 -2422 2500
rect 6822 520 6922 2500
rect -2360 358 6760 458
<< locali >>
rect -2522 2500 -2422 2662
rect -2522 358 -2422 520
rect 6822 2500 6922 2662
rect 6822 358 6922 520
rect 442 -570 490 -562
rect 442 -610 444 -570
rect -2522 -1680 -2422 -1518
rect -2522 -3782 -2422 -3620
rect 6822 -1680 6922 -1518
rect 6822 -3782 6922 -3620
<< viali >>
rect -2422 2562 -2360 2662
rect -2360 2562 6760 2662
rect 6760 2562 6822 2662
rect -2522 563 -2422 2457
rect 6822 563 6922 2457
rect -2422 358 -2360 458
rect -2360 358 6760 458
rect 6760 358 6822 458
rect -1782 -482 -1736 -442
rect 208 -518 256 -470
rect 2674 -490 2714 -450
rect 3274 -530 3308 46
rect 5050 -530 5086 44
rect 5170 -530 5206 44
rect 6172 -530 6208 44
rect 444 -612 492 -570
rect -2044 -714 -1996 -666
rect -320 -716 -272 -668
rect 118 -708 166 -668
rect 352 -710 400 -668
rect 526 -710 574 -668
rect 764 -708 812 -668
rect 1204 -716 1252 -668
rect 2934 -696 2982 -648
rect 676 -828 724 -780
rect 3276 -1208 3310 -852
rect 5052 -1208 5086 -854
rect 5172 -1208 5206 -854
rect 6174 -1208 6208 -852
rect -2422 -1618 -2360 -1518
rect -2360 -1618 6760 -1518
rect 6760 -1618 6822 -1518
rect -2522 -3584 -2422 -1716
rect 6822 -3584 6922 -1716
rect -2422 -3782 -2360 -3682
rect -2360 -3782 6760 -3682
rect 6760 -3782 6822 -3682
<< metal1 >>
rect -2528 2662 6928 2668
rect -2528 2562 -2422 2662
rect 6822 2562 6928 2662
rect -2528 2556 6928 2562
rect -2528 2457 -2416 2556
rect -2528 563 -2522 2457
rect -2422 563 -2416 2457
rect -1816 2256 -1806 2556
rect 6206 2256 6216 2556
rect 6816 2457 6928 2556
rect -2340 2140 6730 2174
rect -2340 2030 -2302 2140
rect 6694 2030 6730 2140
rect -2340 1992 6730 2030
rect -2304 1774 -2298 1834
rect -2238 1774 -2232 1834
rect -2146 1806 -2086 1992
rect -1724 1806 -1664 1992
rect -2298 636 -2238 1774
rect -2146 1746 -1664 1806
rect -1296 1774 -1290 1834
rect -1230 1774 -1224 1834
rect -432 1828 -372 1992
rect 1286 1828 1346 1992
rect 3002 1832 3062 1992
rect 4716 1832 4776 1992
rect -2146 1228 -2086 1746
rect -1724 1642 -1664 1746
rect -1290 1536 -1230 1774
rect -432 1768 1346 1828
rect 2134 1768 2140 1828
rect 2200 1768 2206 1828
rect 3002 1772 4776 1832
rect -1722 1228 -1662 1348
rect -856 1228 -796 1353
rect -2146 1168 -1662 1228
rect -1296 1168 -1290 1228
rect -1230 1168 -1224 1228
rect -862 1168 -856 1228
rect -796 1168 -790 1228
rect -2146 648 -2086 1168
rect -1722 1042 -1662 1168
rect -1290 942 -1230 1168
rect -856 1042 -796 1168
rect -432 946 -372 1768
rect -6 1228 54 1348
rect 426 1228 486 1470
rect 856 1228 916 1350
rect -12 1168 -6 1228
rect 54 1168 60 1228
rect 420 1168 426 1228
rect 486 1168 492 1228
rect 850 1168 856 1228
rect 916 1168 922 1228
rect -6 1050 54 1168
rect 856 1050 916 1168
rect 1286 930 1346 1768
rect 2140 1530 2200 1768
rect 1712 1228 1772 1348
rect 2564 1228 2624 1350
rect 1706 1168 1712 1228
rect 1772 1168 1778 1228
rect 2138 1168 2144 1228
rect 2204 1168 2210 1228
rect 2558 1168 2564 1228
rect 2624 1168 2630 1228
rect 1712 1044 1772 1168
rect 2144 938 2204 1168
rect 2564 1044 2624 1168
rect 3002 934 3062 1772
rect 3426 1228 3486 1348
rect 3860 1228 3920 1470
rect 4296 1228 4356 1346
rect 3420 1168 3426 1228
rect 3486 1168 3492 1228
rect 3854 1168 3860 1228
rect 3920 1168 3926 1228
rect 4290 1168 4296 1228
rect 4356 1168 4362 1228
rect 3426 1048 3486 1168
rect 4296 1048 4356 1168
rect 4716 940 4776 1772
rect 5568 1768 5574 1828
rect 5634 1768 5640 1828
rect 6000 1820 6060 1992
rect 6432 1820 6492 1992
rect 5574 1554 5634 1768
rect 6000 1760 6492 1820
rect 6588 1768 6594 1828
rect 6654 1768 6660 1828
rect 6000 1644 6060 1760
rect 5136 1228 5196 1348
rect 5130 1168 5136 1228
rect 5196 1168 5202 1228
rect 5570 1168 5576 1228
rect 5636 1168 5642 1228
rect 6000 1226 6060 1350
rect 6432 1226 6492 1760
rect 5136 1048 5196 1168
rect 5576 938 5636 1168
rect 6000 1166 6492 1226
rect 6000 1044 6060 1166
rect -1726 648 -1666 748
rect -2304 576 -2298 636
rect -2238 576 -2232 636
rect -2146 588 -1666 648
rect 426 636 486 854
rect 3856 636 3916 858
rect 5996 644 6056 750
rect 6432 644 6492 1166
rect -2528 464 -2416 563
rect -2146 464 -2086 588
rect -1726 464 -1666 588
rect 420 576 426 636
rect 486 576 492 636
rect 3850 576 3856 636
rect 3916 576 3922 636
rect 5996 584 6494 644
rect 6594 636 6654 1768
rect 5996 464 6056 584
rect 6432 464 6492 584
rect 6588 576 6594 636
rect 6654 576 6660 636
rect 6816 563 6822 2457
rect 6922 563 6928 2457
rect 6816 464 6928 563
rect -2528 458 6928 464
rect -2528 358 -2422 458
rect 6822 358 6928 458
rect -2528 352 6928 358
rect -2066 -428 -1822 352
rect -1794 -442 -1728 -370
rect -1066 -428 -822 352
rect -66 -428 178 352
rect 934 -428 1178 352
rect 1934 -428 2178 352
rect 2660 -424 2724 -376
rect -1794 -482 -1782 -442
rect -1736 -482 -1728 -442
rect 2660 -450 2726 -424
rect 2750 -428 2994 352
rect 3260 156 3324 352
rect 3376 156 3436 352
rect 3510 156 3570 352
rect 3634 156 3694 352
rect 3260 96 3694 156
rect 3260 46 3324 96
rect 202 -464 262 -458
rect -1794 -496 -1728 -482
rect 196 -524 202 -464
rect 262 -524 268 -464
rect 2660 -490 2674 -450
rect 2714 -490 2726 -450
rect 2660 -502 2726 -490
rect 202 -530 262 -524
rect 3260 -530 3274 46
rect 3308 -530 3324 46
rect 3376 -72 3436 96
rect 3510 10 3570 96
rect 3634 -94 3694 96
rect 4022 156 4082 352
rect 4152 156 4212 352
rect 4280 156 4340 352
rect 4798 164 4858 352
rect 4928 164 4988 352
rect 4022 96 4340 156
rect 4534 98 4540 158
rect 4600 98 4606 158
rect 4022 10 4082 96
rect 4152 -84 4212 96
rect 4280 8 4340 96
rect 4540 7 4600 98
rect 4662 96 4668 156
rect 4728 96 4734 156
rect 4798 104 4988 164
rect 4668 -96 4728 96
rect 4798 7 4858 104
rect 4928 -107 4988 104
rect 5034 159 5224 352
rect 5274 159 5334 352
rect 5404 159 5464 352
rect 5656 240 5662 300
rect 5722 240 5728 300
rect 5034 99 5464 159
rect 5034 44 5224 99
rect 3260 -540 3324 -530
rect -660 -570 1586 -564
rect -660 -612 444 -570
rect 492 -612 1586 -570
rect 3764 -574 3824 -488
rect 3892 -574 3952 -384
rect -660 -624 1586 -612
rect -2292 -666 -1984 -660
rect -2292 -714 -2044 -666
rect -1996 -714 -1984 -666
rect -2292 -720 -1984 -714
rect -660 -768 -600 -624
rect 436 -626 496 -624
rect 348 -662 408 -656
rect 840 -662 900 -656
rect -332 -668 348 -662
rect -332 -716 -320 -668
rect -272 -708 118 -668
rect 166 -708 348 -668
rect -272 -716 348 -708
rect -332 -722 348 -716
rect 408 -722 412 -662
rect 514 -668 840 -662
rect 514 -710 526 -668
rect 574 -708 764 -668
rect 812 -708 840 -668
rect 574 -710 840 -708
rect 514 -722 840 -710
rect 900 -668 1264 -662
rect 900 -716 1204 -668
rect 1252 -716 1264 -668
rect 900 -722 1264 -716
rect 348 -728 408 -722
rect 840 -728 900 -722
rect 1526 -766 1586 -624
rect 3632 -634 3952 -574
rect 2922 -648 3104 -642
rect 2922 -696 2934 -648
rect 2982 -696 3104 -648
rect 2922 -702 3104 -696
rect 670 -774 730 -768
rect 664 -834 670 -774
rect 730 -834 736 -774
rect 670 -840 730 -834
rect 3262 -852 3326 -840
rect -2066 -1512 -1822 -942
rect -1066 -1512 -822 -942
rect -66 -1512 178 -942
rect 934 -1512 1178 -942
rect 1934 -1512 2178 -942
rect 2752 -1512 2996 -942
rect 3262 -1208 3276 -852
rect 3310 -1208 3326 -852
rect 3632 -982 3692 -634
rect 4410 -744 4470 -398
rect 5034 -530 5050 44
rect 5086 -530 5170 44
rect 5206 -530 5224 44
rect 5274 -98 5334 99
rect 5404 2 5464 99
rect 5526 96 5532 156
rect 5592 96 5598 156
rect 5532 -92 5592 96
rect 5662 -2 5722 240
rect 5920 164 5980 352
rect 6044 164 6104 352
rect 6158 164 6222 352
rect 5920 104 6222 164
rect 5920 2 5980 104
rect 6044 -84 6104 104
rect 6158 44 6222 104
rect 5034 -544 5224 -530
rect 4410 -804 4598 -744
rect 4410 -982 4470 -804
rect 4538 -894 4598 -804
rect 5032 -854 5226 -832
rect 3262 -1258 3326 -1208
rect 3376 -1258 3436 -1072
rect 3510 -1258 3570 -1172
rect 3262 -1318 3570 -1258
rect 3262 -1512 3326 -1318
rect 3376 -1512 3436 -1318
rect 3510 -1512 3570 -1318
rect 3754 -1394 3814 -1172
rect 3748 -1454 3754 -1394
rect 3814 -1454 3820 -1394
rect 3892 -1396 3952 -1086
rect 4022 -1260 4082 -1170
rect 4150 -1260 4210 -1082
rect 4280 -1260 4340 -1172
rect 4022 -1320 4340 -1260
rect 3886 -1456 3892 -1396
rect 3952 -1456 3958 -1396
rect 4022 -1512 4082 -1320
rect 4150 -1512 4210 -1320
rect 4280 -1512 4340 -1320
rect 4666 -1272 4726 -1080
rect 4794 -1272 4854 -1172
rect 4922 -1272 4982 -1080
rect 5032 -1208 5052 -854
rect 5086 -1208 5172 -854
rect 5206 -1208 5226 -854
rect 5788 -970 5848 -406
rect 6158 -530 6172 44
rect 6208 -530 6222 44
rect 6158 -542 6222 -530
rect 6158 -852 6226 -834
rect 5032 -1270 5226 -1208
rect 5274 -1270 5334 -1082
rect 5402 -1270 5462 -1166
rect 5530 -1182 5590 -1088
rect 5530 -1248 5592 -1182
rect 5032 -1272 5462 -1270
rect 4666 -1330 5462 -1272
rect 4666 -1332 5226 -1330
rect 5032 -1512 5226 -1332
rect 5532 -1392 5592 -1248
rect 5666 -1274 5726 -1167
rect 5660 -1334 5666 -1274
rect 5726 -1334 5732 -1274
rect 5916 -1276 5976 -1166
rect 6048 -1276 6108 -1094
rect 6158 -1208 6174 -852
rect 6208 -1208 6226 -852
rect 6158 -1276 6226 -1208
rect 5532 -1458 5592 -1452
rect 5916 -1336 6226 -1276
rect 5916 -1512 5976 -1336
rect 6048 -1512 6108 -1336
rect 6158 -1512 6226 -1336
rect -2528 -1518 6928 -1512
rect -2528 -1618 -2422 -1518
rect 6822 -1618 6928 -1518
rect -2528 -1624 6928 -1618
rect -2528 -1716 -2416 -1624
rect 3892 -1674 3952 -1670
rect 5532 -1674 5592 -1668
rect 3892 -1676 5532 -1674
rect -2528 -3584 -2522 -1716
rect -2422 -3584 -2416 -1716
rect 2526 -1736 3892 -1676
rect 3952 -1734 5532 -1676
rect -1764 -1848 -48 -1788
rect 12 -1848 18 -1788
rect 1664 -1848 1670 -1788
rect 1730 -1848 1736 -1788
rect -1764 -2344 -1704 -1848
rect -1340 -1946 -1280 -1848
rect -48 -2042 12 -1848
rect 1670 -2032 1730 -1848
rect 2526 -2026 2586 -1736
rect 3892 -1742 3952 -1736
rect 5532 -1740 5592 -1734
rect 6816 -1716 6928 -1624
rect 2944 -1848 2950 -1788
rect 3010 -1848 3016 -1788
rect 3382 -1848 3388 -1788
rect 3448 -1848 3454 -1788
rect 5092 -1848 5098 -1788
rect 5158 -1848 6018 -1788
rect 2950 -1948 3010 -1848
rect 3388 -2036 3448 -1848
rect 5098 -2046 5158 -1848
rect 5518 -1946 5578 -1848
rect -1348 -2344 -1288 -2224
rect -908 -2340 -848 -2124
rect -476 -2340 -416 -2224
rect 378 -2340 438 -2218
rect 810 -2340 870 -2134
rect 1230 -2340 1290 -2218
rect 2094 -2340 2154 -2226
rect 3818 -2340 3878 -2226
rect 4244 -2340 4304 -2122
rect 4666 -2340 4726 -2226
rect 5516 -2336 5576 -2222
rect 5958 -2336 6018 -1848
rect -1764 -2404 -1288 -2344
rect -914 -2400 -908 -2340
rect -848 -2400 -842 -2340
rect -482 -2400 -476 -2340
rect -416 -2400 -410 -2340
rect -58 -2400 -52 -2340
rect 8 -2400 14 -2340
rect 372 -2400 378 -2340
rect 438 -2400 444 -2340
rect 804 -2400 810 -2340
rect 870 -2400 876 -2340
rect 1224 -2400 1230 -2340
rect 1290 -2400 1296 -2340
rect 2088 -2400 2094 -2340
rect 2154 -2400 2160 -2340
rect 2944 -2400 2950 -2340
rect 3010 -2400 3016 -2340
rect 3378 -2400 3384 -2340
rect 3444 -2400 3450 -2340
rect 3812 -2400 3818 -2340
rect 3878 -2400 3884 -2340
rect 4238 -2400 4244 -2340
rect 4304 -2400 4310 -2340
rect 4660 -2400 4666 -2340
rect 4726 -2400 4732 -2340
rect 5094 -2400 5100 -2340
rect 5160 -2400 5166 -2340
rect 5516 -2396 6018 -2336
rect -1764 -2892 -1704 -2404
rect -1348 -2526 -1288 -2404
rect -908 -2406 -848 -2400
rect -476 -2530 -416 -2400
rect -52 -2626 8 -2400
rect 378 -2522 438 -2400
rect 2094 -2526 2154 -2400
rect 2950 -2526 3010 -2400
rect 3384 -2636 3444 -2400
rect 3818 -2530 3878 -2400
rect 4666 -2522 4726 -2400
rect 5100 -2618 5160 -2400
rect 5516 -2526 5576 -2396
rect -1340 -2892 -1280 -2800
rect -906 -2892 -846 -2722
rect -1764 -2952 -846 -2892
rect -1764 -3082 -1704 -2952
rect -1340 -3082 -1280 -2952
rect -906 -3082 -846 -2952
rect 808 -2906 868 -2700
rect 1234 -2906 1294 -2804
rect 1670 -2904 1730 -2696
rect 808 -2966 1294 -2906
rect 1664 -2964 1670 -2904
rect 1730 -2964 1736 -2904
rect 808 -3082 868 -2966
rect 1234 -3082 1294 -2966
rect 2526 -3082 2586 -2736
rect 4242 -3082 4302 -2700
rect 5516 -2904 5576 -2800
rect 5958 -2904 6018 -2396
rect 5516 -2964 6018 -2904
rect 5516 -3082 5576 -2964
rect 5958 -3082 6018 -2964
rect -1820 -3122 6120 -3082
rect -1820 -3266 -1782 -3122
rect 6080 -3266 6120 -3122
rect -1820 -3296 6120 -3266
rect -2528 -3676 -2416 -3584
rect -1816 -3676 -1806 -3376
rect 6206 -3676 6216 -3376
rect 6816 -3584 6822 -1716
rect 6922 -3584 6928 -1716
rect 6816 -3676 6928 -3584
rect -2528 -3682 6928 -3676
rect -2528 -3782 -2422 -3682
rect 6822 -3782 6928 -3682
rect -2528 -3788 6928 -3782
<< via1 >>
rect -2416 2256 -1816 2556
rect 6216 2256 6816 2556
rect -2302 2030 6694 2140
rect -2298 1774 -2238 1834
rect -1290 1774 -1230 1834
rect 2140 1768 2200 1828
rect -1290 1168 -1230 1228
rect -856 1168 -796 1228
rect -6 1168 54 1228
rect 426 1168 486 1228
rect 856 1168 916 1228
rect 1712 1168 1772 1228
rect 2144 1168 2204 1228
rect 2564 1168 2624 1228
rect 3426 1168 3486 1228
rect 3860 1168 3920 1228
rect 4296 1168 4356 1228
rect 5574 1768 5634 1828
rect 6594 1768 6654 1828
rect 5136 1168 5196 1228
rect 5576 1168 5636 1228
rect -2298 576 -2238 636
rect 426 576 486 636
rect 3856 576 3916 636
rect 6594 576 6654 636
rect 202 -470 262 -464
rect 202 -518 208 -470
rect 208 -518 256 -470
rect 256 -518 262 -470
rect 202 -524 262 -518
rect 4540 98 4600 158
rect 4668 96 4728 156
rect 5662 240 5722 300
rect 348 -668 408 -662
rect 348 -710 352 -668
rect 352 -710 400 -668
rect 400 -710 408 -668
rect 348 -722 408 -710
rect 840 -722 900 -662
rect 670 -780 730 -774
rect 670 -828 676 -780
rect 676 -828 724 -780
rect 724 -828 730 -780
rect 670 -834 730 -828
rect 5532 96 5592 156
rect 3754 -1454 3814 -1394
rect 3892 -1456 3952 -1396
rect 5666 -1334 5726 -1274
rect 5532 -1452 5592 -1392
rect 3892 -1736 3952 -1676
rect 5532 -1734 5592 -1674
rect -48 -1848 12 -1788
rect 1670 -1848 1730 -1788
rect 2950 -1848 3010 -1788
rect 3388 -1848 3448 -1788
rect 5098 -1848 5158 -1788
rect -908 -2400 -848 -2340
rect -476 -2400 -416 -2340
rect -52 -2400 8 -2340
rect 378 -2400 438 -2340
rect 810 -2400 870 -2340
rect 1230 -2400 1290 -2340
rect 2094 -2400 2154 -2340
rect 2950 -2400 3010 -2340
rect 3384 -2400 3444 -2340
rect 3818 -2400 3878 -2340
rect 4244 -2400 4304 -2340
rect 4666 -2400 4726 -2340
rect 5100 -2400 5160 -2340
rect 1670 -2964 1730 -2904
rect -1782 -3266 6080 -3122
rect -2416 -3676 -1816 -3376
rect 6216 -3676 6816 -3376
<< metal2 >>
rect -2416 2556 -1816 2566
rect -2416 2246 -1816 2256
rect 6216 2556 6816 2566
rect 6216 2246 6816 2256
rect -2340 2140 6730 2174
rect -2340 2030 -2302 2140
rect 6694 2030 6730 2140
rect -2340 1992 6730 2030
rect -2298 1834 -2238 1840
rect -1290 1834 -1230 1840
rect -2238 1774 -1290 1834
rect -2298 1768 -2238 1774
rect -1290 1768 -1230 1774
rect 2140 1828 2200 1834
rect 5574 1828 5634 1834
rect 6594 1828 6654 1834
rect 2200 1768 5574 1828
rect 5634 1768 6594 1828
rect 2140 1762 2200 1768
rect 5574 1762 5634 1768
rect 6594 1762 6654 1768
rect -1290 1228 -1230 1234
rect -856 1228 -796 1234
rect -6 1228 54 1234
rect 426 1228 486 1234
rect 856 1228 916 1234
rect 1712 1228 1772 1234
rect 2144 1228 2204 1234
rect 2564 1228 2624 1234
rect 3426 1228 3486 1234
rect 3860 1228 3920 1234
rect 4296 1228 4356 1234
rect 5136 1228 5196 1234
rect 5576 1228 5636 1234
rect -1230 1168 -856 1228
rect -796 1168 -6 1228
rect 54 1168 426 1228
rect 486 1168 856 1228
rect 916 1168 1712 1228
rect 1772 1168 2144 1228
rect 2204 1168 2564 1228
rect 2624 1168 3426 1228
rect 3486 1168 3860 1228
rect 3920 1168 4296 1228
rect 4356 1168 5136 1228
rect 5196 1168 5576 1228
rect 5636 1168 6776 1228
rect -1290 1162 -1230 1168
rect -856 1162 -796 1168
rect -6 1162 54 1168
rect 426 1162 486 1168
rect 856 1162 916 1168
rect 1712 1162 1772 1168
rect 2144 1162 2204 1168
rect 2564 1162 2624 1168
rect 3426 1162 3486 1168
rect 3860 1162 3920 1168
rect 4296 1162 4356 1168
rect 5136 1162 5196 1168
rect 5576 1162 5636 1168
rect -2298 636 -2238 642
rect 426 636 486 642
rect 3856 636 3916 642
rect 6594 636 6654 642
rect -2238 576 426 636
rect 486 576 3856 636
rect 3916 576 6594 636
rect -2298 570 -2238 576
rect 426 570 486 576
rect 3856 570 3916 576
rect 5662 300 5722 306
rect 202 240 5662 300
rect 202 -464 262 240
rect 5662 234 5722 240
rect 4540 158 4600 164
rect 348 98 4540 158
rect 196 -524 202 -464
rect 262 -524 268 -464
rect 348 -662 408 98
rect 4540 92 4600 98
rect 4668 156 4728 162
rect 5532 156 5592 162
rect 5802 156 5862 576
rect 6594 570 6654 576
rect 4728 96 5532 156
rect 5592 96 5862 156
rect 4668 90 4728 96
rect 5532 90 5592 96
rect 6716 32 6776 1168
rect 6378 -28 6776 32
rect 342 -722 348 -662
rect 408 -722 414 -662
rect 834 -722 840 -662
rect 900 -722 906 -662
rect 664 -834 670 -774
rect 730 -834 736 -774
rect 670 -1394 730 -834
rect 840 -1050 900 -722
rect 840 -1110 3214 -1050
rect 3154 -1274 3214 -1110
rect 5666 -1274 5726 -1268
rect 3154 -1334 5666 -1274
rect 5666 -1340 5726 -1334
rect 3754 -1394 3814 -1388
rect 670 -1454 3754 -1394
rect 3754 -1460 3814 -1454
rect 3892 -1396 3952 -1390
rect 5526 -1452 5532 -1392
rect 5592 -1452 5598 -1392
rect 3892 -1676 3952 -1456
rect 5532 -1674 5592 -1452
rect 3886 -1736 3892 -1676
rect 3952 -1736 3958 -1676
rect 5526 -1734 5532 -1674
rect 5592 -1734 5598 -1674
rect -48 -1788 12 -1782
rect 1670 -1788 1730 -1782
rect 2950 -1788 3010 -1782
rect 3388 -1788 3448 -1782
rect 5098 -1788 5158 -1782
rect 12 -1848 1670 -1788
rect 1730 -1848 2950 -1788
rect 3010 -1848 3388 -1788
rect 3448 -1848 5098 -1788
rect -48 -1854 12 -1848
rect 1670 -1854 1730 -1848
rect 2950 -1854 3010 -1848
rect 3388 -1854 3448 -1848
rect 5098 -1854 5158 -1848
rect -908 -2340 -848 -2334
rect -476 -2340 -416 -2334
rect -52 -2340 8 -2334
rect 378 -2340 438 -2334
rect 810 -2340 870 -2334
rect 1230 -2340 1290 -2334
rect 2094 -2340 2154 -2334
rect 2950 -2340 3010 -2334
rect 3384 -2340 3444 -2334
rect 3818 -2340 3878 -2334
rect 4244 -2340 4304 -2334
rect 4666 -2340 4726 -2334
rect 5100 -2340 5160 -2334
rect -848 -2400 -476 -2340
rect -416 -2400 -52 -2340
rect 8 -2400 378 -2340
rect 438 -2400 810 -2340
rect 870 -2400 1230 -2340
rect 1290 -2400 2094 -2340
rect 2154 -2400 2950 -2340
rect 3010 -2400 3384 -2340
rect 3444 -2400 3818 -2340
rect 3878 -2400 4244 -2340
rect 4304 -2400 4666 -2340
rect 4726 -2400 5100 -2340
rect -908 -2406 -848 -2400
rect -476 -2406 -416 -2400
rect -52 -2406 8 -2400
rect 378 -2406 438 -2400
rect 810 -2406 870 -2400
rect 1230 -2406 1290 -2400
rect 2094 -2406 2154 -2400
rect 2950 -2406 3010 -2400
rect 3384 -2406 3444 -2400
rect 3818 -2406 3878 -2400
rect 4244 -2406 4304 -2400
rect 4666 -2406 4726 -2400
rect 5100 -2406 5160 -2400
rect 1670 -2904 1730 -2898
rect 6378 -2904 6438 -28
rect 1730 -2964 6438 -2904
rect 1670 -2970 1730 -2964
rect -1820 -3122 6120 -3082
rect -1820 -3266 -1782 -3122
rect 6080 -3266 6120 -3122
rect -1820 -3296 6120 -3266
rect -2416 -3376 -1816 -3366
rect -2416 -3686 -1816 -3676
rect 6216 -3376 6816 -3366
rect 6216 -3686 6816 -3676
<< via2 >>
rect -2416 2256 -1816 2556
rect 6216 2256 6816 2556
rect -2302 2030 6694 2140
rect -1782 -3266 6080 -3122
rect -2416 -3676 -1816 -3376
rect 6216 -3676 6816 -3376
<< metal3 >>
rect -2426 2556 -1806 2561
rect -2426 2256 -2416 2556
rect -1816 2256 -1806 2556
rect -2426 2251 -1806 2256
rect 6206 2556 6826 2561
rect 6206 2256 6216 2556
rect 6816 2256 6826 2556
rect 6206 2251 6826 2256
rect -2340 2140 6730 2174
rect -2340 2030 -2302 2140
rect 6694 2030 6730 2140
rect -2340 1992 6730 2030
rect -1820 -3122 6120 -3082
rect -1820 -3266 -1782 -3122
rect 6080 -3266 6120 -3122
rect -1820 -3296 6120 -3266
rect -2426 -3376 -1806 -3371
rect -2426 -3676 -2416 -3376
rect -1816 -3676 -1806 -3376
rect -2426 -3681 -1806 -3676
rect 6206 -3376 6826 -3371
rect 6206 -3676 6216 -3376
rect 6816 -3676 6826 -3376
rect 6206 -3681 6826 -3676
<< via3 >>
rect -2416 2256 -1816 2556
rect 6216 2256 6816 2556
rect -2302 2030 6694 2140
rect -1782 -3266 6080 -3122
rect -2416 -3676 -1816 -3376
rect 6216 -3676 6816 -3376
<< metal4 >>
rect -2600 2556 7000 2740
rect -2600 2256 -2416 2556
rect -1816 2256 6216 2556
rect 6816 2256 7000 2556
rect -2600 2140 7000 2256
rect -2600 2030 -2302 2140
rect 6694 2030 7000 2140
rect -2600 1940 7000 2030
rect -2600 -3122 7000 -3060
rect -2600 -3266 -1782 -3122
rect 6080 -3266 7000 -3122
rect -2600 -3376 7000 -3266
rect -2600 -3676 -2416 -3376
rect -1816 -3676 6216 -3376
rect 6816 -3676 7000 -3376
rect -2600 -3860 7000 -3676
use sky130_fd_pr__nfet_01v8_58Q5WU  sky130_fd_pr__nfet_01v8_58Q5WU_0
timestamp 1623971255
transform 1 0 2128 0 1 -2084
box -3890 -188 3890 188
use sky130_fd_pr__nfet_01v8_58Q5WU  sky130_fd_pr__nfet_01v8_58Q5WU_1
timestamp 1623971255
transform 1 0 2128 0 1 -2666
box -3890 -188 3890 188
use sky130_fd_pr__nfet_01v8_lvt_V7QMZR  sky130_fd_pr__nfet_01v8_lvt_V7QMZR_0
timestamp 1623971255
transform 1 0 5689 0 1 -1031
box -554 -310 554 310
use sky130_fd_pr__nfet_01v8_N6QVV6  sky130_fd_pr__nfet_01v8_N6QVV6_0
timestamp 1623971255
transform 1 0 4180 0 1 -1031
box -941 -310 941 310
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623971255
transform -1 0 604 0 1 -924
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_SCHXZ7  sky130_fd_pr__pfet_01v8_SCHXZ7_0
timestamp 1623971255
transform 1 0 4180 0 1 -244
box -941 -419 941 419
use sky130_fd_pr__pfet_01v8_lvt_HJ2CZP  sky130_fd_pr__pfet_01v8_lvt_HJ2CZP_0
timestamp 1623971255
transform 1 0 5689 0 1 -244
box -554 -419 554 419
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623971255
transform -1 0 880 0 1 -924
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1623971255
transform 1 0 52 0 1 -924
box -38 -48 314 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623375787
transform 1 0 -2064 0 1 -924
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_0
timestamp 1623375787
transform -1 0 2996 0 1 -924
box -38 -48 2154 592
use sky130_fd_pr__pfet_01v8_2Q5KMA  sky130_fd_pr__pfet_01v8_2Q5KMA_1
timestamp 1623971255
transform 1 0 2173 0 1 896
box -4355 -200 4355 200
use sky130_fd_pr__pfet_01v8_2Q5KMA  sky130_fd_pr__pfet_01v8_2Q5KMA_0
timestamp 1623971255
transform 1 0 2173 0 1 1496
box -4355 -200 4355 200
<< labels >>
flabel metal1 2548 -1880 2560 -1874 1 FreeSans 480 0 0 0 vswitchl
flabel metal2 1694 -2378 1704 -2366 1 FreeSans 480 0 0 0 ibiasn
flabel metal1 3656 -862 3666 -854 1 FreeSans 480 0 0 0 vpdiode
flabel metal1 5552 -1226 5564 -1208 1 FreeSans 480 0 0 0 vswitchl
flabel metal2 4962 114 4976 132 1 FreeSans 480 0 0 0 vswitchh
flabel metal2 1104 596 1120 610 1 FreeSans 480 0 0 0 vswitchh
flabel metal1 5812 -840 5822 -830 1 FreeSans 480 0 0 0 vcp
flabel metal1 620 -692 624 -688 1 FreeSans 480 0 0 0 vQB
flabel metal1 294 -700 300 -692 1 FreeSans 480 0 0 0 vQA
flabel metal1 -2200 -692 -2194 -688 1 FreeSans 480 0 0 0 vsig_in
flabel metal1 3070 -680 3078 -676 1 FreeSans 480 0 0 0 vin_div
flabel metal1 300 -592 304 -588 1 FreeSans 480 0 0 0 vRSTN
flabel metal2 944 -1420 952 -1412 1 FreeSans 480 0 0 0 VQBb
flabel metal2 220 -146 228 -138 1 FreeSans 480 0 0 0 vQAb
flabel metal2 1582 1194 1598 1204 1 FreeSans 480 0 0 0 vpbias
flabel metal2 2204 -2944 2214 -2936 1 FreeSans 480 0 0 0 vpbias
flabel metal4 886 2206 898 2222 1 FreeSans 480 0 0 0 VDD
flabel metal4 1252 -3422 1278 -3396 1 FreeSans 480 0 0 0 VSS
flabel metal1 4436 -580 4442 -570 1 FreeSans 480 0 0 0 vndiode
<< properties >>
string FIXED_BBOX -2472 -3732 6872 -1668
<< end >>

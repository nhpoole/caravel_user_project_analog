magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nwell >>
rect -358 582 11058 2438
<< pwell >>
rect -358 -3058 11058 418
<< psubdiff >>
rect -322 282 -160 382
rect 10860 282 11022 382
rect -322 220 -222 282
rect -322 -2922 -222 -2860
rect 10922 220 11022 282
rect 10922 -2922 11022 -2860
rect -322 -3022 -160 -2922
rect 10860 -3022 11022 -2922
<< nsubdiff >>
rect -322 2302 -160 2402
rect 10860 2302 11022 2402
rect -322 2240 -222 2302
rect -322 718 -222 780
rect 10922 2240 11022 2302
rect 10922 718 11022 780
rect -322 618 -160 718
rect 10860 618 11022 718
<< psubdiffcont >>
rect -160 282 10860 382
rect -322 -2860 -222 220
rect 10922 -2860 11022 220
rect -160 -3022 10860 -2922
<< nsubdiffcont >>
rect -160 2302 10860 2402
rect -322 780 -222 2240
rect 10922 780 11022 2240
rect -160 618 10860 718
<< locali >>
rect -322 2242 -222 2402
rect -322 618 -222 778
rect 10922 2242 11022 2402
rect 10922 618 11022 778
rect -322 220 -222 382
rect -322 -3022 -222 -2860
rect 10922 220 11022 382
rect 10922 -3022 11022 -2860
<< viali >>
rect -222 2302 -160 2402
rect -160 2302 10860 2402
rect 10860 2302 10922 2402
rect -322 2240 -222 2242
rect -322 780 -222 2240
rect -322 778 -222 780
rect 10922 2240 11022 2242
rect 10922 780 11022 2240
rect 10922 778 11022 780
rect -222 618 -160 718
rect -160 618 10860 718
rect 10860 618 10922 718
rect -222 282 -160 382
rect -160 282 10860 382
rect 10860 282 10922 382
rect -322 -2762 -222 122
rect 10922 -2762 11022 122
rect -222 -3022 -160 -2922
rect -160 -3022 10860 -2922
rect 10860 -3022 10922 -2922
<< metal1 >>
rect -328 2402 11028 2408
rect -328 2302 -222 2402
rect 10922 2302 11028 2402
rect -328 2296 11028 2302
rect -328 2242 -216 2296
rect -328 778 -322 2242
rect -222 778 -216 2242
rect 384 1996 394 2296
rect 10306 1996 10316 2296
rect 10916 2242 11028 2296
rect 3466 1910 7322 1950
rect 3466 1758 3514 1910
rect 7278 1758 7322 1910
rect 3466 1720 7322 1758
rect -328 724 -216 778
rect 3504 1503 3564 1720
rect 3640 1503 3700 1720
rect 3504 1443 3700 1503
rect 3504 956 3564 1443
rect 3640 1336 3700 1443
rect 4022 1248 4082 1720
rect 4412 1498 4472 1720
rect 4538 1498 4598 1720
rect 4412 1438 4598 1498
rect 4412 1334 4472 1438
rect 3636 956 3696 1042
rect 3504 896 3696 956
rect 3504 724 3564 896
rect 3636 724 3696 896
rect 3764 952 3824 1142
rect 3896 952 3956 1042
rect 4152 952 4212 1042
rect 3764 892 4152 952
rect 4212 892 4218 952
rect 4280 842 4340 1125
rect 4280 776 4340 782
rect 4538 724 4598 1438
rect 4926 1503 4986 1720
rect 5054 1503 5114 1720
rect 5178 1503 5238 1720
rect 5302 1556 5308 1616
rect 5368 1556 5374 1616
rect 4926 1443 5238 1503
rect 4926 1336 4986 1443
rect 4668 952 4728 1042
rect 4662 892 4668 952
rect 4728 892 4734 952
rect 4794 840 4854 1157
rect 4794 774 4854 780
rect 4926 956 4986 1042
rect 5054 956 5114 1443
rect 5178 1332 5238 1443
rect 5308 1238 5368 1556
rect 5568 1248 5628 1720
rect 5958 1497 6018 1720
rect 6086 1497 6146 1720
rect 6218 1497 6278 1720
rect 5958 1437 6278 1497
rect 5958 1334 6018 1437
rect 5182 956 5242 1042
rect 4926 896 5242 956
rect 4926 724 4986 896
rect 5054 724 5114 896
rect 5182 724 5242 896
rect 5440 950 5500 1046
rect 5700 950 5760 1040
rect 5826 950 5886 1140
rect 5440 890 5886 950
rect 5956 950 6016 1044
rect 6086 950 6146 1437
rect 6218 1336 6278 1437
rect 6340 1434 6346 1494
rect 6406 1434 6412 1494
rect 6210 950 6270 1042
rect 5956 890 6270 950
rect 5700 838 5760 890
rect 5700 772 5760 778
rect 5956 724 6016 890
rect 6086 724 6146 890
rect 6210 724 6270 890
rect 6346 948 6406 1434
rect 6472 948 6532 1049
rect 6346 888 6532 948
rect 6602 724 6662 1720
rect 6988 1496 7048 1720
rect 7118 1496 7178 1720
rect 6988 1436 7178 1496
rect 6988 1336 7048 1436
rect 6736 948 6796 1045
rect 6864 948 6924 1148
rect 6736 888 6924 948
rect 6864 836 6924 888
rect 6988 952 7048 1044
rect 7118 952 7178 1436
rect 6988 892 7178 952
rect 6858 776 6864 836
rect 6924 776 6930 836
rect 6988 724 7048 892
rect 7118 724 7178 892
rect 10916 778 10922 2242
rect 11022 778 11028 2242
rect 10916 724 11028 778
rect -328 718 11028 724
rect -328 618 -222 718
rect 10922 618 11028 718
rect -328 612 11028 618
rect 3052 524 3112 530
rect 5700 524 5760 530
rect 8088 524 8148 530
rect 3112 464 5700 524
rect 5760 464 8088 524
rect 3052 458 3112 464
rect 5700 458 5760 464
rect 8088 458 8148 464
rect -328 382 11028 388
rect -328 282 -222 382
rect 10922 282 11028 382
rect -328 276 11028 282
rect -328 122 -216 276
rect -328 -2762 -322 122
rect -222 4 -216 122
rect 726 4 786 276
rect 852 4 912 276
rect 1488 170 1494 230
rect 1554 170 1560 230
rect 2524 170 2530 230
rect 2590 170 2596 230
rect 974 54 980 114
rect 1040 54 1046 114
rect -222 -56 912 4
rect -222 -728 -216 -56
rect 726 -728 786 -56
rect 852 -140 912 -56
rect 980 -240 1040 54
rect 1364 -56 1370 4
rect 1430 -56 1436 4
rect 1370 -146 1430 -56
rect 1494 -236 1554 170
rect 2006 54 2012 114
rect 2072 54 2078 114
rect 1618 -56 1624 4
rect 1684 -56 1690 4
rect 1624 -142 1684 -56
rect 2012 -250 2072 54
rect 2390 -56 2396 4
rect 2456 -56 2462 4
rect 2396 -150 2456 -56
rect 2530 -240 2590 170
rect 3042 54 3048 114
rect 3108 54 3114 114
rect 2652 -56 2658 4
rect 2718 -56 2724 4
rect 2658 -142 2718 -56
rect 3048 -246 3108 54
rect 3172 4 3232 276
rect 3306 4 3366 276
rect 4022 4 4082 276
rect 4146 4 4206 276
rect 4784 176 4790 236
rect 4850 176 4856 236
rect 5820 176 5826 236
rect 5886 176 5892 236
rect 4270 60 4276 120
rect 4336 60 4342 120
rect 3172 -56 4206 4
rect 3172 -138 3232 -56
rect 852 -728 912 -622
rect 1110 -726 1170 -618
rect -222 -788 912 -728
rect 1104 -786 1110 -726
rect 1170 -786 1176 -726
rect -222 -2762 -216 -788
rect 26 -896 32 -836
rect 92 -896 98 -836
rect 32 -2170 92 -896
rect 172 -1082 232 -788
rect 1240 -836 1300 -546
rect 1752 -836 1812 -546
rect 1886 -726 1946 -622
rect 2140 -726 2200 -620
rect 1880 -786 1886 -726
rect 1946 -786 1952 -726
rect 2134 -786 2140 -726
rect 2200 -786 2206 -726
rect 2272 -836 2332 -542
rect 2788 -836 2848 -542
rect 2918 -726 2978 -622
rect 2912 -786 2918 -726
rect 2978 -786 2984 -726
rect 3172 -728 3232 -616
rect 3306 -728 3366 -56
rect 4022 -728 4082 -56
rect 4146 -144 4206 -56
rect 4276 -234 4336 60
rect 4660 -50 4666 10
rect 4726 -50 4732 10
rect 4666 -140 4726 -50
rect 4790 -230 4850 176
rect 5302 60 5308 120
rect 5368 60 5374 120
rect 4914 -50 4920 10
rect 4980 -50 4986 10
rect 4920 -136 4980 -50
rect 5308 -244 5368 60
rect 5686 -50 5692 10
rect 5752 -50 5758 10
rect 5692 -144 5752 -50
rect 5826 -234 5886 176
rect 6338 60 6344 120
rect 6404 60 6410 120
rect 5948 -50 5954 10
rect 6014 -50 6020 10
rect 5954 -136 6014 -50
rect 6344 -240 6404 60
rect 6470 10 6530 276
rect 6602 10 6662 276
rect 7318 10 7378 276
rect 7442 10 7502 276
rect 8080 170 8086 230
rect 8146 170 8152 230
rect 9116 170 9122 230
rect 9182 170 9188 230
rect 7566 54 7572 114
rect 7632 54 7638 114
rect 6470 -50 7502 10
rect 6470 -144 6530 -50
rect 4148 -728 4208 -616
rect 4406 -720 4466 -612
rect 1746 -896 1752 -836
rect 1812 -896 1818 -836
rect 2266 -896 2272 -836
rect 2332 -896 2338 -836
rect 2782 -896 2788 -836
rect 2848 -896 2854 -836
rect 1240 -902 1300 -896
rect 2918 -958 2978 -786
rect 3172 -788 4208 -728
rect 4400 -780 4406 -720
rect 4466 -780 4472 -720
rect 2912 -1018 2918 -958
rect 2978 -1018 2984 -958
rect 172 -1142 654 -1082
rect 1024 -1142 1030 -1082
rect 1090 -1142 1096 -1082
rect 172 -1632 232 -1142
rect 594 -1246 654 -1142
rect 1030 -1336 1090 -1142
rect 596 -1632 656 -1524
rect 1456 -1626 1516 -1524
rect 172 -1692 656 -1632
rect 1026 -1686 1032 -1626
rect 1092 -1686 1516 -1626
rect 172 -2162 232 -1692
rect 596 -1792 656 -1692
rect 1032 -1890 1092 -1686
rect 1456 -1786 1516 -1686
rect 592 -2162 652 -2070
rect 26 -2230 32 -2170
rect 92 -2230 98 -2170
rect 172 -2222 652 -2162
rect 172 -2336 232 -2222
rect 592 -2336 652 -2222
rect 1890 -2336 1950 -1394
rect 2314 -1626 2374 -1520
rect 2748 -1626 2808 -1424
rect 3178 -1626 3238 -1520
rect 2308 -1682 2314 -1626
rect 2374 -1682 2380 -1626
rect 2308 -1686 2380 -1682
rect 2742 -1686 2748 -1626
rect 2808 -1686 2814 -1626
rect 2314 -1788 2374 -1686
rect 2748 -1866 2808 -1686
rect 3178 -1788 3238 -1682
rect 3606 -2336 3666 -788
rect 4536 -830 4596 -540
rect 4536 -1082 4596 -890
rect 4798 -958 4858 -478
rect 5048 -830 5108 -540
rect 5182 -720 5242 -616
rect 5436 -720 5496 -614
rect 5176 -780 5182 -720
rect 5242 -780 5248 -720
rect 5430 -780 5436 -720
rect 5496 -780 5502 -720
rect 5568 -830 5628 -536
rect 6084 -830 6144 -536
rect 6214 -720 6274 -616
rect 6208 -780 6214 -720
rect 6274 -780 6280 -720
rect 6468 -722 6528 -610
rect 6602 -722 6662 -50
rect 7318 -722 7378 -50
rect 7442 -140 7502 -50
rect 7572 -240 7632 54
rect 7956 -56 7962 4
rect 8022 -56 8028 4
rect 7962 -146 8022 -56
rect 8086 -236 8146 170
rect 8598 54 8604 114
rect 8664 54 8670 114
rect 8210 -56 8216 4
rect 8276 -56 8282 4
rect 8216 -142 8276 -56
rect 8604 -250 8664 54
rect 8982 -56 8988 4
rect 9048 -56 9054 4
rect 8988 -150 9048 -56
rect 9122 -240 9182 170
rect 9634 54 9640 114
rect 9700 54 9706 114
rect 9244 -56 9250 4
rect 9310 -56 9316 4
rect 9250 -142 9310 -56
rect 9640 -246 9700 54
rect 9766 2 9826 276
rect 9898 2 9958 276
rect 10916 122 11028 276
rect 10916 2 10922 122
rect 9766 -58 10922 2
rect 9766 -140 9826 -58
rect 7444 -722 7504 -618
rect 6468 -782 7504 -722
rect 7702 -726 7762 -618
rect 5042 -890 5048 -830
rect 5108 -890 5114 -830
rect 5562 -890 5568 -830
rect 5628 -890 5634 -830
rect 6078 -890 6084 -830
rect 6144 -890 6150 -830
rect 4792 -1018 4798 -958
rect 4858 -1018 4864 -958
rect 4458 -1142 4464 -1082
rect 4524 -1142 4596 -1082
rect 4894 -1140 5818 -1080
rect 4464 -1340 4524 -1142
rect 4894 -1248 4954 -1140
rect 4038 -1626 4098 -1520
rect 4896 -1624 4956 -1520
rect 5320 -1624 5380 -1140
rect 5758 -1248 5818 -1140
rect 5756 -1624 5816 -1520
rect 4038 -1788 4098 -1682
rect 4462 -1686 4468 -1626
rect 4528 -1686 4534 -1626
rect 4896 -1684 5816 -1624
rect 6184 -1626 6244 -1426
rect 6610 -1626 6670 -1520
rect 4468 -1890 4528 -1686
rect 4896 -1788 4956 -1684
rect 4894 -2168 4954 -2064
rect 5320 -2168 5380 -1684
rect 5756 -1788 5816 -1684
rect 6178 -1686 6184 -1626
rect 6244 -1686 6250 -1626
rect 6604 -1682 6610 -1626
rect 6670 -1682 6676 -1626
rect 6604 -1686 6676 -1682
rect 6610 -1788 6670 -1686
rect 5756 -2168 5816 -2062
rect 4894 -2228 5816 -2168
rect 6180 -2170 6240 -1984
rect 4894 -2336 4954 -2228
rect 5320 -2336 5380 -2228
rect 5756 -2336 5816 -2228
rect 6174 -2230 6180 -2170
rect 6240 -2230 6246 -2170
rect 7038 -2336 7098 -782
rect 7696 -786 7702 -726
rect 7762 -786 7768 -726
rect 7832 -836 7892 -546
rect 8344 -836 8404 -546
rect 8478 -726 8538 -622
rect 8732 -726 8792 -620
rect 8472 -786 8478 -726
rect 8538 -786 8544 -726
rect 8726 -786 8732 -726
rect 8792 -786 8798 -726
rect 8864 -836 8924 -542
rect 9380 -836 9440 -542
rect 9510 -726 9570 -622
rect 9504 -786 9510 -726
rect 9570 -786 9576 -726
rect 9764 -728 9824 -616
rect 9898 -728 9958 -58
rect 10916 -728 10922 -58
rect 9764 -788 10922 -728
rect 7826 -896 7832 -836
rect 7892 -896 7898 -836
rect 8338 -896 8344 -836
rect 8404 -896 8410 -836
rect 8858 -896 8864 -836
rect 8924 -896 8930 -836
rect 9374 -896 9380 -836
rect 9440 -896 9446 -836
rect 9608 -1026 9614 -966
rect 9674 -1026 9680 -966
rect 9614 -1332 9674 -1026
rect 10044 -1096 10104 -788
rect 10468 -1096 10528 -788
rect 10594 -896 10600 -836
rect 10660 -896 10666 -836
rect 10044 -1156 10528 -1096
rect 10044 -1246 10104 -1156
rect 7468 -1626 7528 -1520
rect 7896 -1626 7956 -1410
rect 8322 -1626 8382 -1520
rect 7468 -1788 7528 -1682
rect 7890 -1686 7896 -1626
rect 7956 -1686 7962 -1626
rect 7896 -1880 7956 -1686
rect 8322 -1788 8382 -1682
rect 8756 -2336 8816 -1418
rect 9186 -1620 9246 -1520
rect 9186 -1626 9248 -1620
rect 9186 -1686 9188 -1626
rect 9186 -1692 9248 -1686
rect 10042 -1630 10102 -1520
rect 10468 -1630 10528 -1156
rect 10042 -1690 10528 -1630
rect 9186 -1788 9246 -1692
rect 10042 -1788 10102 -1690
rect 9612 -2164 9672 -1982
rect 10044 -2164 10104 -2066
rect 10468 -2164 10528 -1690
rect 10600 -2164 10660 -896
rect 9606 -2224 9612 -2164
rect 9672 -2224 9678 -2164
rect 10044 -2224 10528 -2164
rect 10594 -2224 10600 -2164
rect 10660 -2224 10666 -2164
rect 10044 -2336 10104 -2224
rect 10468 -2336 10528 -2224
rect -66 -2384 10708 -2336
rect -66 -2494 -4 -2384
rect 10652 -2494 10708 -2384
rect -66 -2550 10708 -2494
rect -328 -2916 -216 -2762
rect 384 -2916 394 -2616
rect 10306 -2916 10316 -2616
rect 10916 -2762 10922 -788
rect 11022 -2762 11028 122
rect 10916 -2916 11028 -2762
rect -328 -2922 11028 -2916
rect -328 -3022 -222 -2922
rect 10922 -3022 11028 -2922
rect -328 -3028 11028 -3022
<< via1 >>
rect -216 1996 384 2296
rect 10316 1996 10916 2296
rect 3514 1758 7278 1910
rect 4152 892 4212 952
rect 4280 782 4340 842
rect 5308 1556 5368 1616
rect 4668 892 4728 952
rect 4794 780 4854 840
rect 6346 1434 6406 1494
rect 5700 778 5760 838
rect 6864 776 6924 836
rect 3052 464 3112 524
rect 5700 464 5760 524
rect 8088 464 8148 524
rect 1494 170 1554 230
rect 2530 170 2590 230
rect 980 54 1040 114
rect 1370 -56 1430 4
rect 2012 54 2072 114
rect 1624 -56 1684 4
rect 2396 -56 2456 4
rect 3048 54 3108 114
rect 2658 -56 2718 4
rect 4790 176 4850 236
rect 5826 176 5886 236
rect 4276 60 4336 120
rect 1110 -786 1170 -726
rect 32 -896 92 -836
rect 1886 -786 1946 -726
rect 2140 -786 2200 -726
rect 2918 -786 2978 -726
rect 4666 -50 4726 10
rect 5308 60 5368 120
rect 4920 -50 4980 10
rect 5692 -50 5752 10
rect 6344 60 6404 120
rect 5954 -50 6014 10
rect 8086 170 8146 230
rect 9122 170 9182 230
rect 7572 54 7632 114
rect 1240 -896 1300 -836
rect 1752 -896 1812 -836
rect 2272 -896 2332 -836
rect 2788 -896 2848 -836
rect 4406 -780 4466 -720
rect 2918 -1018 2978 -958
rect 1030 -1142 1090 -1082
rect 1032 -1686 1092 -1626
rect 32 -2230 92 -2170
rect 2314 -1682 2374 -1626
rect 2748 -1686 2808 -1626
rect 3178 -1682 3238 -1626
rect 4536 -890 4596 -830
rect 5182 -780 5242 -720
rect 5436 -780 5496 -720
rect 6214 -780 6274 -720
rect 7962 -56 8022 4
rect 8604 54 8664 114
rect 8216 -56 8276 4
rect 8988 -56 9048 4
rect 9640 54 9700 114
rect 9250 -56 9310 4
rect 5048 -890 5108 -830
rect 5568 -890 5628 -830
rect 6084 -890 6144 -830
rect 4798 -1018 4858 -958
rect 4464 -1142 4524 -1082
rect 4038 -1682 4098 -1626
rect 4468 -1686 4528 -1626
rect 6184 -1686 6244 -1626
rect 6610 -1682 6670 -1626
rect 6180 -2230 6240 -2170
rect 7702 -786 7762 -726
rect 8478 -786 8538 -726
rect 8732 -786 8792 -726
rect 9510 -786 9570 -726
rect 7832 -896 7892 -836
rect 8344 -896 8404 -836
rect 8864 -896 8924 -836
rect 9380 -896 9440 -836
rect 9614 -1026 9674 -966
rect 10600 -896 10660 -836
rect 7468 -1682 7528 -1626
rect 7896 -1686 7956 -1626
rect 8322 -1682 8382 -1626
rect 9188 -1686 9248 -1626
rect 9612 -2224 9672 -2164
rect 10600 -2224 10660 -2164
rect -4 -2494 10652 -2384
rect -216 -2916 384 -2616
rect 10316 -2916 10916 -2616
<< metal2 >>
rect -216 2296 384 2306
rect -216 1986 384 1996
rect 10316 2296 10916 2306
rect 10316 1986 10916 1996
rect 3466 1910 7322 1950
rect 3466 1758 3514 1910
rect 7278 1758 7322 1910
rect 3466 1720 7322 1758
rect 5308 1616 5368 1622
rect 602 1556 5308 1616
rect 602 168 662 1556
rect 5308 1550 5368 1556
rect 6346 1494 6406 1500
rect 2532 1434 6346 1494
rect 2532 236 2592 1434
rect 6346 1428 6406 1434
rect 4152 952 4212 958
rect 4668 952 4728 958
rect 4212 892 4668 952
rect 4728 892 10792 952
rect 4152 886 4212 892
rect 4668 886 4728 892
rect 4274 782 4280 842
rect 4340 782 4346 842
rect 3046 464 3052 524
rect 3112 464 3118 524
rect -84 108 662 168
rect 1494 230 1554 236
rect 2530 230 2592 236
rect 1554 170 2530 230
rect 2590 170 2592 230
rect 1494 164 1554 170
rect 2530 164 2590 170
rect 3052 120 3112 464
rect 4280 126 4340 782
rect 4788 780 4794 840
rect 4854 780 4860 840
rect 4794 242 4854 780
rect 5694 778 5700 838
rect 5760 778 5766 838
rect 6864 836 6924 842
rect 5700 524 5760 778
rect 6924 776 7632 836
rect 6864 770 6924 776
rect 5694 464 5700 524
rect 5760 464 5766 524
rect 4790 236 4854 242
rect 5826 236 5886 242
rect 4850 176 5826 236
rect 4790 170 4850 176
rect 5826 170 5886 176
rect 980 114 1040 120
rect 2012 114 2072 120
rect 3048 114 3112 120
rect -84 -1626 -24 108
rect 1040 54 2012 114
rect 2072 54 3048 114
rect 3108 54 3112 114
rect 4276 120 4340 126
rect 5308 120 5368 126
rect 6344 120 6404 126
rect 4336 60 5308 120
rect 5368 60 6344 120
rect 6404 60 7262 120
rect 4276 54 4336 60
rect 5308 54 5368 60
rect 6344 54 6404 60
rect 980 48 1040 54
rect 2012 48 2072 54
rect 3048 48 3108 54
rect 4666 10 4726 16
rect 4920 10 4980 16
rect 5692 10 5752 16
rect 5954 10 6014 16
rect 1370 4 1430 10
rect 1624 4 1684 10
rect 2396 4 2456 10
rect 2658 4 2718 10
rect 1430 -56 1624 4
rect 1684 -56 2396 4
rect 2456 -56 2658 4
rect 2718 -56 3716 4
rect 4726 -50 4920 10
rect 4980 -50 5692 10
rect 5752 -50 5954 10
rect 4666 -56 4726 -50
rect 4920 -56 4980 -50
rect 5692 -56 5752 -50
rect 5954 -56 6014 -50
rect 7202 4 7262 60
rect 7572 114 7632 776
rect 8082 464 8088 524
rect 8148 464 8154 524
rect 8088 236 8148 464
rect 8086 230 8148 236
rect 9122 230 9182 236
rect 8146 170 9122 230
rect 8086 164 8146 170
rect 9122 164 9182 170
rect 8604 114 8664 120
rect 9640 114 9700 120
rect 7632 54 8604 114
rect 8664 54 9640 114
rect 7572 48 7632 54
rect 8604 48 8664 54
rect 9640 48 9700 54
rect 7962 4 8022 10
rect 8216 4 8276 10
rect 8988 4 9048 10
rect 9250 4 9310 10
rect 7202 -56 7962 4
rect 8022 -56 8216 4
rect 8276 -56 8988 4
rect 9048 -56 9250 4
rect 1370 -62 1430 -56
rect 1624 -62 1684 -56
rect 2396 -62 2456 -56
rect 2658 -62 2718 -56
rect 1110 -726 1170 -720
rect 1886 -726 1946 -720
rect 2140 -726 2200 -720
rect 2918 -726 2978 -720
rect 1170 -786 1886 -726
rect 1946 -786 2140 -726
rect 2200 -786 2918 -726
rect 1110 -792 1170 -786
rect 1886 -792 1946 -786
rect 2140 -792 2200 -786
rect 2918 -792 2978 -786
rect 32 -836 92 -830
rect 1752 -836 1812 -830
rect 2272 -836 2332 -830
rect 2788 -836 2848 -830
rect 92 -896 1240 -836
rect 1300 -896 1752 -836
rect 1812 -896 2272 -836
rect 2332 -896 2788 -836
rect 3656 -838 3716 -56
rect 7962 -62 8022 -56
rect 8216 -62 8276 -56
rect 8988 -62 9048 -56
rect 9250 -62 9310 -56
rect 4406 -720 4466 -714
rect 5182 -720 5242 -714
rect 5436 -720 5496 -714
rect 6214 -720 6274 -714
rect 4466 -780 5182 -720
rect 5242 -780 5436 -720
rect 5496 -780 6214 -720
rect 4406 -786 4466 -780
rect 5182 -786 5242 -780
rect 5436 -786 5496 -780
rect 6214 -786 6274 -780
rect 7702 -726 7762 -720
rect 8478 -726 8538 -720
rect 8732 -726 8792 -720
rect 9510 -726 9570 -720
rect 7762 -786 8478 -726
rect 8538 -786 8732 -726
rect 8792 -786 9510 -726
rect 7702 -792 7764 -786
rect 8478 -792 8538 -786
rect 8732 -792 8792 -786
rect 9510 -792 9570 -786
rect 5048 -830 5108 -824
rect 5568 -830 5628 -824
rect 6084 -830 6144 -824
rect 32 -902 92 -896
rect 1752 -902 1812 -896
rect 2272 -902 2332 -896
rect 2788 -902 2848 -896
rect 3647 -898 3656 -838
rect 3716 -898 3725 -838
rect 4530 -890 4536 -830
rect 4596 -890 5048 -830
rect 5108 -890 5568 -830
rect 5628 -890 6084 -830
rect 7704 -840 7764 -792
rect 7832 -836 7892 -830
rect 8344 -836 8404 -830
rect 8864 -836 8924 -830
rect 9380 -836 9440 -830
rect 10600 -836 10660 -830
rect 5048 -896 5108 -890
rect 5568 -896 5628 -890
rect 6084 -896 6144 -890
rect 7697 -896 7706 -840
rect 7762 -896 7771 -840
rect 7892 -896 8344 -836
rect 8404 -896 8864 -836
rect 8924 -896 9380 -836
rect 9440 -896 10600 -836
rect 7704 -898 7764 -896
rect 7832 -902 7892 -896
rect 8344 -902 8404 -896
rect 8864 -902 8924 -896
rect 9380 -902 9440 -896
rect 10600 -902 10660 -896
rect 2918 -958 2978 -952
rect 4798 -958 4858 -952
rect 2978 -1018 4798 -958
rect 2918 -1024 2978 -1018
rect 4798 -1024 4858 -1018
rect 9614 -966 9674 -960
rect 10732 -966 10792 892
rect 9674 -1026 10792 -966
rect 9614 -1032 9674 -1026
rect 1030 -1082 1090 -1076
rect 4464 -1082 4524 -1076
rect 1090 -1142 4464 -1082
rect 1030 -1148 1090 -1142
rect 4464 -1148 4524 -1142
rect 1032 -1626 1092 -1620
rect -84 -1686 1032 -1626
rect 1032 -1692 1092 -1686
rect 2314 -1626 2374 -1620
rect 2748 -1626 2808 -1620
rect 4468 -1626 4528 -1620
rect 6184 -1626 6244 -1620
rect 6610 -1626 6670 -1620
rect 7896 -1626 7956 -1620
rect 2374 -1682 2748 -1626
rect 2314 -1686 2748 -1682
rect 2808 -1682 3178 -1626
rect 3238 -1682 4038 -1626
rect 4098 -1682 4468 -1626
rect 2808 -1686 4468 -1682
rect 4528 -1686 6184 -1626
rect 6244 -1682 6610 -1626
rect 6670 -1682 7468 -1626
rect 7528 -1682 7896 -1626
rect 6244 -1686 7896 -1682
rect 7956 -1682 8322 -1626
rect 8382 -1682 9188 -1626
rect 7956 -1686 9188 -1682
rect 9248 -1686 9254 -1626
rect 2314 -1692 2374 -1686
rect 2748 -1692 2808 -1686
rect 4468 -1692 4528 -1686
rect 6184 -1692 6244 -1686
rect 6610 -1692 6670 -1686
rect 7896 -1692 7956 -1686
rect 9612 -2164 9672 -2158
rect 10600 -2164 10660 -2158
rect 32 -2170 92 -2164
rect 6180 -2170 6240 -2164
rect 92 -2230 6180 -2170
rect 9672 -2224 10600 -2164
rect 9612 -2230 9672 -2224
rect 10600 -2230 10660 -2224
rect 32 -2236 92 -2230
rect 6180 -2236 6240 -2230
rect -66 -2384 10708 -2336
rect -66 -2494 -4 -2384
rect 10652 -2494 10708 -2384
rect -66 -2550 10708 -2494
rect -216 -2616 384 -2606
rect -216 -2926 384 -2916
rect 10316 -2616 10916 -2606
rect 10316 -2926 10916 -2916
<< via2 >>
rect -216 1996 384 2296
rect 10316 1996 10916 2296
rect 3514 1758 7278 1910
rect 3656 -898 3716 -838
rect 7706 -896 7762 -840
rect -4 -2494 10652 -2384
rect -216 -2916 384 -2616
rect 10316 -2916 10916 -2616
<< metal3 >>
rect -226 2296 394 2301
rect -226 1996 -216 2296
rect 384 1996 394 2296
rect -226 1991 394 1996
rect 10306 2296 10926 2301
rect 10306 1996 10316 2296
rect 10916 1996 10926 2296
rect 10306 1991 10926 1996
rect 3466 1910 7322 1950
rect 3466 1758 3514 1910
rect 7278 1758 7322 1910
rect 3466 1720 7322 1758
rect 3628 -838 7786 -820
rect 3628 -898 3656 -838
rect 3716 -840 7786 -838
rect 3716 -896 7706 -840
rect 7762 -896 7786 -840
rect 3716 -898 7786 -896
rect 3628 -920 7786 -898
rect -66 -2384 10708 -2336
rect -66 -2494 -4 -2384
rect 10652 -2494 10708 -2384
rect -66 -2550 10708 -2494
rect -226 -2616 394 -2611
rect -226 -2916 -216 -2616
rect 384 -2916 394 -2616
rect -226 -2921 394 -2916
rect 10306 -2616 10926 -2611
rect 10306 -2916 10316 -2616
rect 10916 -2916 10926 -2616
rect 10306 -2921 10926 -2916
<< via3 >>
rect -216 1996 384 2296
rect 10316 1996 10916 2296
rect 3514 1758 7278 1910
rect -4 -2494 10652 -2384
rect -216 -2916 384 -2616
rect 10316 -2916 10916 -2616
<< metal4 >>
rect -400 2296 11100 2480
rect -400 1996 -216 2296
rect 384 1996 10316 2296
rect 10916 1996 11100 2296
rect -400 1910 11100 1996
rect -400 1758 3514 1910
rect 7278 1758 11100 1910
rect -400 1680 11100 1758
rect -400 -2384 11100 -2300
rect -400 -2494 -4 -2384
rect 10652 -2494 11100 -2384
rect -400 -2616 11100 -2494
rect -400 -2916 -216 -2616
rect 384 -2916 10316 -2616
rect 10916 -2916 11100 -2616
rect -400 -3100 11100 -2916
use sky130_fd_pr__nfet_01v8_YXNJ6N  sky130_fd_pr__nfet_01v8_YXNJ6N_1
timestamp 1623971255
transform 1 0 8635 0 1 -378
box -1319 -288 1319 288
use sky130_fd_pr__nfet_01v8_3YN2WN  sky130_fd_pr__nfet_01v8_3YN2WN_0
timestamp 1623971255
transform 1 0 5353 0 1 -1386
box -5177 -188 5177 188
use sky130_fd_pr__nfet_01v8_3YN2WN  sky130_fd_pr__nfet_01v8_3YN2WN_1
timestamp 1623971255
transform 1 0 5353 0 1 -1926
box -5177 -188 5177 188
use sky130_fd_pr__pfet_01v8_HVERXA  sky130_fd_pr__pfet_01v8_HVERXA_0
timestamp 1623971255
transform 1 0 5343 0 1 1190
box -1871 -200 1871 200
use sky130_fd_pr__nfet_01v8_lvt_YXNJ6N  sky130_fd_pr__nfet_01v8_lvt_YXNJ6N_0
timestamp 1623971255
transform 1 0 5339 0 1 -378
box -1319 -288 1319 288
use sky130_fd_pr__nfet_01v8_YXNJ6N  sky130_fd_pr__nfet_01v8_YXNJ6N_0
timestamp 1623971255
transform 1 0 2043 0 1 -378
box -1319 -288 1319 288
<< labels >>
flabel metal1 1044 -1164 1062 -1152 1 FreeSans 480 0 0 0 vtail_diff
flabel metal1 9634 -1132 9650 -1116 1 FreeSans 480 0 0 0 vbiasp
flabel metal1 9628 -2132 9644 -2122 1 FreeSans 480 0 0 0 vcmn_tail2
flabel metal1 6202 -2146 6214 -2134 1 FreeSans 480 0 0 0 vcmn_tail1
flabel metal1 1262 -1662 1270 -1654 1 FreeSans 480 0 0 0 vcmc
flabel metal2 6878 -1662 6892 -1652 1 FreeSans 480 0 0 0 ibiasn
flabel metal2 8640 -872 8650 -858 1 FreeSans 480 0 0 0 vcmn_tail2
flabel metal2 8428 -30 8440 -14 1 FreeSans 480 0 0 0 vom
flabel metal2 8082 -768 8104 -750 1 FreeSans 480 0 0 0 vocm
flabel metal2 7816 84 7828 94 1 FreeSans 480 0 0 0 vcmcn2
flabel metal2 8638 196 8648 208 1 FreeSans 480 0 0 0 vcmcn
flabel metal2 4368 918 4374 930 1 FreeSans 480 0 0 0 vbiasp
flabel metal2 5334 -876 5352 -860 1 FreeSans 480 0 0 0 vtail_diff
flabel metal2 5154 -28 5172 -12 1 FreeSans 480 0 0 0 vim
flabel metal2 4486 84 4506 96 1 FreeSans 480 0 0 0 vom
flabel metal2 5310 198 5330 214 1 FreeSans 480 0 0 0 vop
flabel metal2 2032 190 2050 210 1 FreeSans 480 0 0 0 vcmcn1
flabel metal2 1136 72 1156 86 1 FreeSans 480 0 0 0 vcmcn
flabel metal2 1856 -42 1878 -30 1 FreeSans 480 0 0 0 vocm
flabel metal2 1492 -760 1510 -748 1 FreeSans 480 0 0 0 vop
flabel metal2 2030 -874 2050 -858 1 FreeSans 480 0 0 0 vcmn_tail1
flabel metal2 4684 -754 4692 -748 1 FreeSans 480 0 0 0 vip
flabel metal1 5328 1322 5346 1338 1 FreeSans 480 0 0 0 vcmc
flabel metal2 4306 554 4312 558 1 FreeSans 480 0 0 0 vom
flabel metal2 4818 552 4824 558 1 FreeSans 480 0 0 0 vop
flabel metal4 -66 2456 -54 2470 1 FreeSans 480 0 0 0 VDD
flabel metal4 172 -3088 186 -3074 1 FreeSans 480 0 0 0 VSS
<< properties >>
string FIXED_BBOX -272 -2972 10972 332
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623986634
<< metal1 >>
rect 23080 14160 23140 14166
rect 23140 14100 24468 14160
rect 23080 14094 23140 14100
rect 27146 14096 27152 14196
rect 27252 14096 27258 14196
rect 32380 14118 32930 14178
rect 29948 8646 30222 8706
<< via1 >>
rect 23080 14100 23140 14160
rect 27152 14096 27252 14196
<< metal2 >>
rect 27152 14196 27252 14202
rect 23074 14100 23080 14160
rect 23140 14100 23146 14160
rect 27148 14101 27152 14191
rect 27252 14101 27256 14191
rect 23080 9432 23140 14100
rect 27152 14090 27252 14096
rect 34621 13582 34630 13642
rect 34690 13582 34699 13642
rect 30988 12438 32238 12498
rect 34630 8592 34690 13582
<< via2 >>
rect 27157 14101 27247 14191
rect 34630 13582 34690 13642
<< metal3 >>
rect 27152 14191 27252 14196
rect 27152 14101 27157 14191
rect 27247 14101 27252 14191
rect 27152 13664 27252 14101
rect 27152 13642 34698 13664
rect 27152 13582 34630 13642
rect 34690 13582 34698 13642
rect 27152 13564 34698 13582
<< metal4 >>
rect 32818 17542 38736 17578
rect 32818 16812 37972 17542
rect 38702 16812 38736 17542
rect 32818 16778 38736 16812
rect 23256 10806 32856 11076
rect 30394 8472 30514 10240
rect 35772 8584 35892 10308
rect 33074 5166 33194 6154
<< via4 >>
rect 37972 16812 38702 17542
<< metal5 >>
rect 37936 17542 38736 17578
rect 37936 16812 37972 17542
rect 38702 16812 38736 17542
rect 37936 6956 38736 16812
use freq_div  freq_div_0 freq_div
timestamp 1623986634
transform 1 0 32794 0 1 8554
box -2674 -2906 3321 454
use cs_ring_osc  cs_ring_osc_0 cs_ring_osc
timestamp 1623971255
transform 1 0 -2466 0 1 6424
box 9760 -28686 41209 4472
use pfd_cp_lpf  pfd_cp_lpf_0 pfd_cp_lpf
timestamp 1623984492
transform -1 0 30256 0 1 14838
box -2600 -3860 7000 2740
<< labels >>
flabel metal1 32888 14140 32900 14154 1 FreeSans 480 0 0 0 vsigin
flabel metal2 32196 12456 32208 12470 1 FreeSans 480 0 0 0 ibiasn
flabel metal4 30452 9650 30462 9664 1 FreeSans 480 0 0 0 VSS
flabel metal4 33486 17114 33506 17132 1 FreeSans 480 0 0 0 VDD
flabel metal1 23198 14118 23210 14134 1 FreeSans 480 0 0 0 vcp
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< metal3 >>
rect -350 -900 244 900
<< mimcap >>
rect -250 760 150 800
rect -250 -760 -210 760
rect 110 -760 150 760
rect -250 -800 150 -760
<< mimcapcontact >>
rect -210 -760 110 760
<< metal4 >>
rect -211 760 111 761
rect -211 -760 -210 760
rect 110 -760 111 760
rect -211 -761 111 -760
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -350 -900 250 900
string parameters w 2.00 l 8.00 val 35.8 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< metal3 >>
rect -1350 -300 1232 300
<< mimcap >>
rect -1250 160 1150 200
rect -1250 -160 -1210 160
rect 1110 -160 1150 160
rect -1250 -200 1150 -160
<< mimcapcontact >>
rect -1210 -160 1110 160
<< metal4 >>
rect -1211 160 1111 161
rect -1211 -160 -1210 160
rect 1110 -160 1111 160
rect -1211 -161 1111 -160
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -1350 -300 1250 300
string parameters w 12.00 l 2.00 val 53.32 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< metal3 >>
rect -350 1272 349 1300
rect -350 -1272 265 1272
rect 329 -1272 349 1272
rect -350 -1300 349 -1272
<< via3 >>
rect 265 -1272 329 1272
<< mimcap >>
rect -250 1160 150 1200
rect -250 -1160 -210 1160
rect 110 -1160 150 1160
rect -250 -1200 150 -1160
<< mimcapcontact >>
rect -210 -1160 110 1160
<< metal4 >>
rect 249 1272 345 1288
rect -211 1160 111 1161
rect -211 -1160 -210 1160
rect 110 -1160 111 1160
rect -211 -1161 111 -1160
rect 249 -1272 265 1272
rect 329 -1272 345 1272
rect 249 -1288 345 -1272
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -350 -1300 250 1300
string parameters w 2.00 l 12.00 val 53.32 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
string library sky130
<< end >>

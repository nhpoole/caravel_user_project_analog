magic
tech sky130A
magscale 1 2
timestamp 1624477805
<< error_s >>
rect 29134 530602 29220 530630
rect 29350 530566 29378 530650
rect 102490 530568 102518 530650
rect 175906 530560 175934 530650
rect 249230 530562 249258 530650
rect 322646 530560 322674 530650
rect 395970 530562 395998 530650
rect 469386 530564 469414 530650
rect 542618 530566 542646 530650
rect 542772 530602 542862 530630
rect 29134 500410 29214 500438
rect 29134 470218 29214 470246
rect 29134 440026 29214 440054
rect 29134 409902 29214 409930
rect 29134 379710 29214 379738
rect 29134 349518 29214 349546
rect 29134 319394 29214 319422
rect 29134 289202 29214 289230
rect 542778 274174 542862 274202
rect 29134 259010 29212 259038
rect 29134 228818 29220 228846
rect 29134 198694 29214 198722
rect 29134 168502 29212 168530
rect 29134 138310 29210 138338
rect 29134 108186 29216 108214
rect 29134 77994 29214 78022
rect 29134 47802 29220 47830
rect 29134 17678 29230 17706
rect 542780 17678 542862 17706
<< nwell >>
rect 97364 586526 98856 587312
<< pwell >>
rect 251660 555238 252036 555720
<< metal1 >>
rect 171904 702112 172024 702118
rect 171904 701868 172024 701992
rect 174410 702112 174530 702118
rect 174410 701868 174530 701992
rect 223692 702112 223812 702118
rect 223692 701868 223812 701992
rect 226092 702112 226212 702118
rect 226092 701868 226212 701992
rect 325330 702112 325450 702118
rect 325330 701868 325450 701992
rect 327840 702112 327960 702118
rect 327840 701868 327960 701992
rect 171904 701150 172024 701262
rect 171904 701024 172024 701030
rect 174410 701150 174530 701262
rect 174410 701024 174530 701030
rect 223692 701150 223812 701262
rect 223692 701024 223812 701030
rect 226092 701150 226212 701262
rect 226092 701024 226212 701030
rect 325330 701150 325450 701262
rect 325330 701024 325450 701030
rect 327840 701150 327960 701262
rect 327840 701024 327960 701030
rect 281522 638598 281582 638604
rect 281050 638538 281522 638598
rect 281522 638532 281582 638538
rect 270574 595388 270674 595394
rect 271642 595388 271742 595394
rect 270674 595288 271642 595388
rect 270574 595282 270674 595288
rect 271642 595282 271742 595288
rect 251483 554476 251773 554522
rect 579046 14540 579052 14662
rect 579174 14542 579299 14662
rect 579899 14542 580143 14662
rect 579174 14540 579267 14542
rect 579928 14540 580143 14542
rect 580265 14540 580271 14662
rect 579058 9814 579064 9936
rect 579186 9816 579311 9936
rect 579911 9816 580155 9936
rect 579186 9814 579279 9816
rect 579940 9814 580155 9816
rect 580277 9814 580283 9936
rect 579170 5084 579176 5206
rect 579298 5084 579391 5206
rect 580052 5084 580267 5206
rect 580389 5084 580395 5206
<< via1 >>
rect 171904 701992 172024 702112
rect 174410 701992 174530 702112
rect 223692 701992 223812 702112
rect 226092 701992 226212 702112
rect 325330 701992 325450 702112
rect 327840 701992 327960 702112
rect 171904 701030 172024 701150
rect 174410 701030 174530 701150
rect 223692 701030 223812 701150
rect 226092 701030 226212 701150
rect 325330 701030 325450 701150
rect 327840 701030 327960 701150
rect 281522 638538 281582 638598
rect 270574 595288 270674 595388
rect 271642 595288 271742 595388
rect 579052 14540 579174 14662
rect 580143 14540 580265 14662
rect 579064 9814 579186 9936
rect 580155 9814 580277 9936
rect 579176 5084 579298 5206
rect 580267 5084 580389 5206
<< metal2 >>
rect 171904 702112 172024 702121
rect 174410 702112 174530 702121
rect 223692 702112 223812 702121
rect 226092 702112 226212 702121
rect 325330 702112 325450 702121
rect 327840 702112 327960 702121
rect 171898 701992 171904 702112
rect 172024 701992 172030 702112
rect 174404 701992 174410 702112
rect 174530 701992 174536 702112
rect 223686 701992 223692 702112
rect 223812 701992 223818 702112
rect 226086 701992 226092 702112
rect 226212 701992 226218 702112
rect 325324 701992 325330 702112
rect 325450 701992 325456 702112
rect 327834 701992 327840 702112
rect 327960 701992 327966 702112
rect 171904 701983 172024 701992
rect 174410 701983 174530 701992
rect 223692 701983 223812 701992
rect 226092 701983 226212 701992
rect 325330 701983 325450 701992
rect 327840 701983 327960 701992
rect 128656 701378 134915 701804
rect 26120 700682 26580 700691
rect 24004 700222 26120 700682
rect 26120 700213 26580 700222
rect 69181 700256 73612 700674
rect 18310 697685 18730 697689
rect 18305 697680 20597 697685
rect 18305 697260 18310 697680
rect 18730 697260 20597 697680
rect 28697 697645 29117 697649
rect 18305 697255 20597 697260
rect 24191 697640 29122 697645
rect 18310 697251 18730 697255
rect 24191 697220 28697 697640
rect 29117 697220 29122 697640
rect 24191 697215 29122 697220
rect 28697 697211 29117 697215
rect 12317 694278 30193 694688
rect 30603 694278 30612 694688
rect 7656 685550 9732 685950
rect 10132 685550 10141 685950
rect 10111 683066 11033 683071
rect 2919 682855 3223 682859
rect 2914 682850 4271 682855
rect 2914 682546 2919 682850
rect 3223 682546 4271 682850
rect 2914 682541 4271 682546
rect 2919 682537 3223 682541
rect 7828 682498 11033 683066
rect 9010 679966 9410 679975
rect 7544 679570 9010 679962
rect 9010 679557 9410 679566
rect 10111 678139 11033 682498
rect 12317 679971 12727 694278
rect 69181 690581 69599 700256
rect 133170 699258 133538 699267
rect 130731 698878 131181 698882
rect 129100 698873 131186 698878
rect 122377 698862 122827 698866
rect 122372 698857 125904 698862
rect 122372 698407 122377 698857
rect 122827 698407 125904 698857
rect 129100 698423 130731 698873
rect 131181 698423 131186 698873
rect 129100 698418 131186 698423
rect 130731 698414 131181 698418
rect 122372 698402 125904 698407
rect 122377 698398 122827 698402
rect 70569 697684 70947 697688
rect 70564 697679 73834 697684
rect 70564 697301 70569 697679
rect 70947 697301 73834 697679
rect 70564 697296 73834 697301
rect 77192 697662 79362 697668
rect 77192 697653 79367 697662
rect 70569 697292 70947 697296
rect 77192 697280 78989 697653
rect 78989 697266 79367 697275
rect 81976 695439 81985 695845
rect 82391 695439 82400 695845
rect 133170 695774 133538 698890
rect 81985 694670 82391 695439
rect 122457 695406 122466 695774
rect 122834 695406 133538 695774
rect 71588 694264 71597 694670
rect 72003 694264 82391 694670
rect 69181 690154 69599 690163
rect 134489 690591 134915 701378
rect 171898 701030 171904 701150
rect 172024 701030 172030 701150
rect 174404 701030 174410 701150
rect 174530 701030 174536 701150
rect 223686 701030 223692 701150
rect 223812 701030 223818 701150
rect 226086 701030 226092 701150
rect 226212 701030 226218 701150
rect 325324 701030 325330 701150
rect 325450 701030 325456 701150
rect 327834 701030 327840 701150
rect 327960 701030 327966 701150
rect 171904 699140 172024 701030
rect 174410 700926 174530 701030
rect 223692 700926 223812 701030
rect 226092 700926 226212 701030
rect 325330 700926 325450 701030
rect 171895 699020 171904 699140
rect 172024 699020 172033 699140
rect 174410 699134 174514 700926
rect 196531 700255 196540 700837
rect 197122 700255 197131 700837
rect 219622 700323 220106 700328
rect 174410 699021 174514 699030
rect 194103 697430 194112 697890
rect 194572 697430 194581 697890
rect 186408 695448 186788 695500
rect 186399 695068 186408 695448
rect 186788 695068 186797 695448
rect 185235 694488 185244 694632
rect 185388 694488 185397 694632
rect 134489 690156 134915 690165
rect 12308 679561 12317 679971
rect 12727 679561 12736 679971
rect 7576 677217 11033 678139
rect 4122 657477 5114 657482
rect 4118 656495 4127 657477
rect 5109 656495 5118 657477
rect 4122 338749 5114 656495
rect 7576 549435 8498 677217
rect 9587 658559 9596 659461
rect 10498 658559 10507 659461
rect 7576 549131 7866 549435
rect 8170 549131 8498 549435
rect 7576 549052 8498 549131
rect 9596 600659 10498 658559
rect 11758 655201 12658 655206
rect 11754 654311 11763 655201
rect 12653 654311 12662 655201
rect 9596 600461 9895 600659
rect 10093 600461 10498 600659
rect 4122 338647 4603 338749
rect 4705 338647 5114 338749
rect 4122 338630 5114 338647
rect 6634 548715 7768 548794
rect 6634 548373 7079 548715
rect 7421 548373 7768 548715
rect 6634 81661 7768 548373
rect 9596 547559 10498 600461
rect 9596 547309 9963 547559
rect 10213 547309 10498 547559
rect 9596 121337 10498 547309
rect 11758 381971 12658 654311
rect 91824 638532 94332 638644
rect 90749 622136 90758 622152
rect 90570 622108 90758 622136
rect 90749 622092 90758 622108
rect 90818 622092 90827 622152
rect 90665 619960 90674 619976
rect 90574 619932 90674 619960
rect 90665 619916 90674 619932
rect 90734 619916 90743 619976
rect 90953 617716 90962 617732
rect 90574 617688 90962 617716
rect 90953 617672 90962 617688
rect 91022 617672 91031 617732
rect 90751 615472 90760 615488
rect 90570 615444 90760 615472
rect 90751 615428 90760 615444
rect 90820 615428 90829 615488
rect 90741 613228 90750 613244
rect 90574 613200 90750 613228
rect 90741 613184 90750 613200
rect 90810 613184 90819 613244
rect 90699 611052 90708 611068
rect 90572 611024 90708 611052
rect 90699 611008 90708 611024
rect 90768 611008 90777 611068
rect 90723 608808 90732 608824
rect 90574 608780 90732 608808
rect 90723 608764 90732 608780
rect 90792 608764 90801 608824
rect 90657 606564 90666 606580
rect 90572 606536 90666 606564
rect 90657 606520 90666 606536
rect 90726 606520 90735 606580
rect 90691 604320 90700 604336
rect 90570 604292 90700 604320
rect 90691 604276 90700 604292
rect 90760 604276 90769 604336
rect 74050 602048 74542 602076
rect 11758 381869 12237 381971
rect 12339 381869 12658 381971
rect 11758 381792 12658 381869
rect 14310 601359 14978 601382
rect 14310 601153 14575 601359
rect 14781 601153 14978 601359
rect 14310 550261 14978 601153
rect 14310 550011 14573 550261
rect 14823 550011 14978 550261
rect 14310 248959 14978 550011
rect 16692 596965 17468 596986
rect 16692 596625 16898 596965
rect 17238 596625 17468 596965
rect 16692 468415 17468 596625
rect 74050 594561 74167 602048
rect 74718 601282 74746 602076
rect 74693 601222 74702 601282
rect 74762 601222 74771 601282
rect 82538 600586 82566 602082
rect 90358 601720 90386 602162
rect 91824 602118 91936 638532
rect 98678 620000 98798 620009
rect 98365 617777 98483 617786
rect 98061 615521 98179 615530
rect 97757 613263 97875 613272
rect 97467 611055 97585 611064
rect 97187 608857 97305 608866
rect 96883 606601 97001 606610
rect 90738 602076 91936 602118
rect 90570 602048 91936 602076
rect 90738 602006 91936 602048
rect 82513 600526 82522 600586
rect 82582 600526 82591 600586
rect 74050 594435 74167 594444
rect 90315 585709 90430 601720
rect 91824 596852 91936 602006
rect 91824 596731 91936 596740
rect 96629 604367 96747 604376
rect 96629 594258 96747 604249
rect 96625 594150 96634 594258
rect 96742 594150 96751 594258
rect 96629 594145 96747 594150
rect 96883 593962 97001 606483
rect 96879 593854 96888 593962
rect 96996 593854 97005 593962
rect 96883 593849 97001 593854
rect 97187 593694 97305 608739
rect 97183 593586 97192 593694
rect 97300 593586 97309 593694
rect 97187 593581 97305 593586
rect 97467 593424 97585 610937
rect 97463 593316 97472 593424
rect 97580 593316 97589 593424
rect 97467 593311 97585 593316
rect 97757 593112 97875 613145
rect 97753 593004 97762 593112
rect 97870 593004 97879 593112
rect 97757 592999 97875 593004
rect 98061 592822 98179 615403
rect 98057 592714 98066 592822
rect 98174 592714 98183 592822
rect 98061 592709 98179 592714
rect 98365 592532 98483 617659
rect 98361 592424 98370 592532
rect 98478 592424 98487 592532
rect 98365 592419 98483 592424
rect 98678 592263 98798 619880
rect 185244 617687 185388 694488
rect 185649 693166 185658 693302
rect 185794 693166 185803 693302
rect 185244 617597 185271 617687
rect 185361 617597 185388 617687
rect 185244 617570 185388 617597
rect 185658 617673 185794 693166
rect 186408 617739 186788 695068
rect 194112 633070 194572 697430
rect 196540 689907 197122 700255
rect 219618 699849 219627 700323
rect 220101 699849 220110 700323
rect 209714 698010 213770 698398
rect 209714 693983 210102 698010
rect 219622 695486 220106 699849
rect 210649 695448 211019 695452
rect 210644 695443 213252 695448
rect 210644 695073 210649 695443
rect 211019 695073 213252 695443
rect 210644 695068 213252 695073
rect 210649 695064 211019 695068
rect 217014 695002 220106 695486
rect 221404 699256 221768 699265
rect 223696 699148 223800 700926
rect 226094 699168 226198 700926
rect 321254 700815 321929 700820
rect 313064 700809 313742 700814
rect 264679 700300 264688 700484
rect 264872 700300 264881 700484
rect 226094 699055 226198 699064
rect 223696 699035 223800 699044
rect 202378 693974 210102 693983
rect 202378 693593 209714 693974
rect 202378 692802 202768 693593
rect 209714 693577 210102 693586
rect 201658 692412 202768 692802
rect 204962 692393 205298 692397
rect 204957 692388 214309 692393
rect 221404 692392 221768 698892
rect 204957 692052 204962 692388
rect 205298 692052 214309 692388
rect 204957 692047 214309 692052
rect 204962 692043 205298 692047
rect 216576 692028 221768 692392
rect 196540 689325 198199 689907
rect 201703 689341 203819 689923
rect 201328 686458 202461 686804
rect 202807 686458 202816 686804
rect 203237 684908 203819 689341
rect 196540 684326 203819 684908
rect 196540 643266 197122 684326
rect 264688 659432 264872 700300
rect 313060 700141 313069 700809
rect 313737 700141 313746 700809
rect 321250 700150 321259 700815
rect 321924 700150 321933 700815
rect 310798 698891 310807 699253
rect 311169 698891 311178 699253
rect 310807 692004 311169 698891
rect 313064 695177 313742 700141
rect 314732 698040 315200 698049
rect 315200 697572 316514 698040
rect 314732 697563 315200 697572
rect 313064 694499 316479 695177
rect 321254 695160 321929 700150
rect 325346 699108 325450 700926
rect 327840 700926 327960 701030
rect 327840 699120 327944 700926
rect 327840 699007 327944 699016
rect 401679 699560 406962 699946
rect 325346 698995 325450 699004
rect 323703 696231 323712 697045
rect 324526 696231 324535 697045
rect 319471 694485 321929 695160
rect 310807 691642 316624 692004
rect 282148 663213 282157 663367
rect 282311 663213 282320 663367
rect 279750 661640 279759 661700
rect 279819 661640 279828 661700
rect 264688 659248 265668 659432
rect 215174 656787 215183 657025
rect 215421 656787 215430 657025
rect 196540 643206 199146 643266
rect 196540 643204 197122 643206
rect 215183 638231 215421 656787
rect 215877 654524 215886 654776
rect 216138 654524 216147 654776
rect 215886 638864 216138 654524
rect 222630 648426 222758 648435
rect 222758 648298 222870 648426
rect 222630 648289 222758 648298
rect 265484 639622 265668 659248
rect 279759 657346 279819 661640
rect 282157 646930 282311 663213
rect 281522 646776 282311 646930
rect 265484 639438 266472 639622
rect 220299 638864 220389 638868
rect 215886 638859 220394 638864
rect 215886 638769 220299 638859
rect 220389 638769 220394 638859
rect 215886 638764 220394 638769
rect 220299 638760 220389 638764
rect 215183 637993 216470 638231
rect 216232 634334 216470 637993
rect 220155 634334 220245 634338
rect 216232 634329 220250 634334
rect 216232 634239 220155 634329
rect 220245 634239 220250 634329
rect 216232 634234 220250 634239
rect 216232 634233 216470 634234
rect 220155 634230 220245 634234
rect 194112 632610 202278 633070
rect 201818 631492 202278 632610
rect 201818 631432 203356 631492
rect 201818 631430 202278 631432
rect 266288 629562 266472 639438
rect 281522 638598 281582 646776
rect 294194 640050 294492 640110
rect 294552 640050 294561 640110
rect 281516 638538 281522 638598
rect 281582 638538 281588 638598
rect 285231 634098 285433 634103
rect 285227 633906 285236 634098
rect 285428 633906 285437 634098
rect 267168 632565 267177 632767
rect 267379 632565 267388 632767
rect 265750 629378 266472 629562
rect 244663 628506 244672 628690
rect 244856 628506 244865 628690
rect 265750 628686 265934 629378
rect 244672 624544 244856 628506
rect 265741 628502 265750 628686
rect 265934 628502 265943 628686
rect 245661 628155 245670 628357
rect 245872 628155 245881 628357
rect 267177 628352 267379 632565
rect 285231 632479 285433 633906
rect 285222 632277 285231 632479
rect 285433 632277 285442 632479
rect 282607 631830 282616 631930
rect 282716 631830 282725 631930
rect 289032 631925 289132 631930
rect 289028 631835 289037 631925
rect 289127 631835 289136 631925
rect 289032 630778 289132 631835
rect 289032 630776 295028 630778
rect 289032 630678 295332 630776
rect 294048 630001 294304 630006
rect 294044 629755 294053 630001
rect 294299 629755 294308 630001
rect 291971 629376 291980 629476
rect 292080 629376 292089 629476
rect 267173 628160 267182 628352
rect 267374 628160 267383 628352
rect 267177 628155 267379 628160
rect 245670 625741 245872 628155
rect 291980 626835 292080 629376
rect 291976 626745 291985 626835
rect 292075 626745 292084 626835
rect 291980 626740 292080 626745
rect 294048 625760 294304 629755
rect 294822 627029 295332 630678
rect 294813 626519 294822 627029
rect 295332 626519 295341 627029
rect 245670 625651 245715 625741
rect 245805 625651 245872 625741
rect 245670 625644 245872 625651
rect 294039 625504 294048 625760
rect 294304 625504 294313 625760
rect 292225 623746 292315 623750
rect 292220 623741 294316 623746
rect 292220 623651 292225 623741
rect 292315 623651 294316 623741
rect 292220 623646 294316 623651
rect 294416 623646 294425 623746
rect 292225 623642 292315 623646
rect 185658 617583 185681 617673
rect 185771 617583 185794 617673
rect 185658 617560 185794 617583
rect 186404 617369 186413 617739
rect 186783 617369 186792 617739
rect 186408 617364 186788 617369
rect 182719 615814 182728 615914
rect 182828 615814 182837 615914
rect 182728 605699 182828 615814
rect 183057 615408 183066 615508
rect 183166 615408 183175 615508
rect 183066 607683 183166 615408
rect 183062 607593 183071 607683
rect 183161 607593 183170 607683
rect 183066 607588 183166 607593
rect 182724 605609 182733 605699
rect 182823 605609 182832 605699
rect 182728 605604 182828 605609
rect 270579 595388 270669 595392
rect 271642 595388 271742 602430
rect 270568 595288 270574 595388
rect 270674 595288 270680 595388
rect 271636 595288 271642 595388
rect 271742 595288 271748 595388
rect 270579 595284 270669 595288
rect 98674 592153 98683 592263
rect 98793 592153 98802 592263
rect 98678 592148 98798 592153
rect 90315 585619 90325 585709
rect 90415 585619 90430 585709
rect 90315 578416 90430 585619
rect 91840 587526 94346 587638
rect 90313 578311 90322 578416
rect 90427 578311 90436 578416
rect 90315 578299 90430 578311
rect 90681 568610 90690 568626
rect 90590 568582 90690 568610
rect 90681 568566 90690 568582
rect 90750 568566 90759 568626
rect 90969 566366 90978 566382
rect 90590 566338 90978 566366
rect 90969 566322 90978 566338
rect 91038 566322 91047 566382
rect 90767 564122 90776 564138
rect 90586 564094 90776 564122
rect 90767 564078 90776 564094
rect 90836 564078 90845 564138
rect 90757 561878 90766 561894
rect 90590 561850 90766 561878
rect 90757 561834 90766 561850
rect 90826 561834 90835 561894
rect 90715 559702 90724 559718
rect 90588 559674 90724 559702
rect 90715 559658 90724 559674
rect 90784 559658 90793 559718
rect 90739 557458 90748 557474
rect 90590 557430 90748 557458
rect 90739 557414 90748 557430
rect 90808 557414 90817 557474
rect 90673 555214 90682 555230
rect 90588 555186 90682 555214
rect 90673 555170 90682 555186
rect 90742 555170 90751 555230
rect 90707 552970 90716 552986
rect 90586 552942 90716 552970
rect 90707 552926 90716 552942
rect 90776 552926 90785 552986
rect 91840 550768 91952 587526
rect 93691 578306 93700 578421
rect 93815 578306 93824 578421
rect 74319 550726 74430 550768
rect 90754 550726 91952 550768
rect 74319 550698 74548 550726
rect 16692 468313 17053 468415
rect 17155 468313 17468 468415
rect 16692 468220 17468 468313
rect 22226 544249 23022 544294
rect 22226 543995 22543 544249
rect 22797 543995 23022 544249
rect 22226 425193 23022 543995
rect 29318 541799 29423 541808
rect 29312 541694 29318 541794
rect 29312 541685 29423 541694
rect 22226 425091 22621 425193
rect 22723 425091 23022 425193
rect 22226 425028 23022 425091
rect 26112 539501 27404 539534
rect 26112 539055 26511 539501
rect 26957 539055 27404 539501
rect 26112 295527 27404 539055
rect 29312 534306 29416 541685
rect 29303 534202 29312 534306
rect 29416 534202 29425 534306
rect 29312 530722 29416 534202
rect 74319 533180 74430 550698
rect 74734 550170 74762 550716
rect 74709 550110 74718 550170
rect 74778 550110 74787 550170
rect 82554 547470 82582 550718
rect 90374 550580 90402 550722
rect 90586 550698 91952 550726
rect 90754 550656 91952 550698
rect 82529 547410 82538 547470
rect 82598 547410 82607 547470
rect 90331 541804 90446 550580
rect 91840 544184 91952 550656
rect 91831 544072 91840 544184
rect 91952 544072 91961 544184
rect 90322 541689 90331 541804
rect 90446 541689 90455 541804
rect 93700 541799 93815 578306
rect 101784 568102 101940 568111
rect 101363 566441 101521 566459
rect 100896 564194 101060 564203
rect 100463 561929 100593 561938
rect 99970 559724 100090 559733
rect 99470 557504 99598 557513
rect 99053 555269 99187 555278
rect 98621 553023 98755 553032
rect 93696 541694 93705 541799
rect 93810 541694 93819 541799
rect 93700 541689 93815 541694
rect 74319 533060 74430 533069
rect 98621 532934 98755 552889
rect 98617 532810 98626 532934
rect 98750 532810 98759 532934
rect 98621 532805 98755 532810
rect 99053 532684 99187 555135
rect 99049 532560 99058 532684
rect 99182 532560 99191 532684
rect 99053 532555 99187 532560
rect 99470 532437 99598 557376
rect 99466 532319 99475 532437
rect 99593 532319 99602 532437
rect 99470 532314 99598 532319
rect 99970 532215 100090 559604
rect 99966 532105 99975 532215
rect 100085 532105 100094 532215
rect 99970 532100 100090 532105
rect 100463 531960 100593 561799
rect 100459 531840 100468 531960
rect 100588 531840 100597 531960
rect 100463 531835 100593 531840
rect 100896 531685 101060 564030
rect 100892 531531 100901 531685
rect 101055 531531 101064 531685
rect 100896 531526 101060 531531
rect 101363 531350 101521 566283
rect 101359 531202 101368 531350
rect 101516 531202 101525 531350
rect 101363 531197 101521 531202
rect 101784 531035 101940 567946
rect 183928 561633 184028 561638
rect 183924 561543 183933 561633
rect 184023 561543 184032 561633
rect 149940 556673 150040 556678
rect 149936 556583 149945 556673
rect 150035 556583 150044 556673
rect 149540 554689 149640 554694
rect 149536 554599 149545 554689
rect 149635 554599 149644 554689
rect 149540 549362 149640 554599
rect 149531 549262 149540 549362
rect 149640 549262 149649 549362
rect 149940 548618 150040 556583
rect 183928 555004 184028 561543
rect 251836 557534 251896 557543
rect 251896 557474 252104 557534
rect 251836 557465 251896 557474
rect 226886 555249 227082 555254
rect 226882 555063 226891 555249
rect 227077 555063 227086 555249
rect 182912 554904 184028 555004
rect 182912 551026 183012 554904
rect 182903 550926 182912 551026
rect 183012 550926 183021 551026
rect 149931 548518 149940 548618
rect 150040 548518 150049 548618
rect 225796 548612 225916 554692
rect 226886 552466 227082 555063
rect 226877 552270 226886 552466
rect 227082 552270 227091 552466
rect 323712 551127 324526 696231
rect 326095 692323 326104 693573
rect 327354 692323 327363 693573
rect 323712 550819 323930 551127
rect 324238 550819 324526 551127
rect 323712 550808 324526 550819
rect 326104 548775 327354 692323
rect 401679 691099 402065 699560
rect 417389 699249 417731 699258
rect 403319 697045 404123 697049
rect 414474 697045 415278 697049
rect 403314 697040 407485 697045
rect 403314 696236 403319 697040
rect 404123 696236 407485 697040
rect 403314 696231 407485 696236
rect 410401 697040 415283 697045
rect 410401 696236 414474 697040
rect 415278 696236 415283 697040
rect 410401 696231 415283 696236
rect 403319 696227 404123 696231
rect 414474 696227 415278 696231
rect 417389 693910 417731 698907
rect 470545 699255 470899 699264
rect 459850 696214 460194 696223
rect 460194 695870 461858 696214
rect 459850 695861 460194 695870
rect 410642 693568 417731 693910
rect 467602 693328 468170 693337
rect 456947 692760 456956 693328
rect 457524 692760 461852 693328
rect 465516 692760 467602 693328
rect 467602 692751 468170 692760
rect 401679 690622 402065 690713
rect 470545 690222 470899 698901
rect 562827 695304 562836 695684
rect 563216 695304 574538 695684
rect 569177 692878 569871 692882
rect 567686 692873 569876 692878
rect 562085 692860 562779 692864
rect 562080 692855 564634 692860
rect 562080 692161 562085 692855
rect 562779 692161 564634 692855
rect 567686 692179 569177 692873
rect 569871 692179 569876 692873
rect 567686 692174 569876 692179
rect 569177 692170 569871 692174
rect 562080 692156 564634 692161
rect 562085 692152 562779 692156
rect 465608 689868 470899 690222
rect 560028 689712 560392 689721
rect 560392 689348 571046 689712
rect 560028 689339 560392 689348
rect 333289 683126 333298 683830
rect 334002 683126 334011 683830
rect 333298 632147 334002 683126
rect 570682 677644 571046 689348
rect 574158 683606 574538 695304
rect 574158 683226 575776 683606
rect 572977 680148 572986 680716
rect 573554 680148 575276 680716
rect 578940 680148 580556 680716
rect 581124 680148 581133 680716
rect 570682 677280 575342 677644
rect 567378 663569 567972 663581
rect 567378 662985 567394 663569
rect 567978 662985 567987 663569
rect 545434 633699 546234 633704
rect 545430 632909 545439 633699
rect 546229 632909 546238 633699
rect 333294 631453 333303 632147
rect 333997 631453 334006 632147
rect 333298 631448 334002 631453
rect 332399 627024 332909 627029
rect 332395 626524 332404 627024
rect 332904 626524 332913 627024
rect 330324 625953 331056 625958
rect 330320 625231 330329 625953
rect 331051 625231 331060 625953
rect 330324 618022 331056 625231
rect 330315 617290 330324 618022
rect 331056 617290 331065 618022
rect 332399 613019 332909 626524
rect 332390 612509 332399 613019
rect 332909 612509 332918 613019
rect 545434 582800 546234 632909
rect 545434 581991 546234 582000
rect 225787 548492 225796 548612
rect 225916 548492 225925 548612
rect 326104 548281 326375 548775
rect 326869 548281 327354 548775
rect 326104 548212 327354 548281
rect 102435 547371 102444 547501
rect 102574 547371 102583 547501
rect 101780 530889 101789 531035
rect 101935 530889 101944 531035
rect 102444 530990 102574 547371
rect 395919 536843 395928 536957
rect 396042 536843 396051 536957
rect 322595 535759 322604 535901
rect 322746 535759 322755 535901
rect 249181 534653 249190 534771
rect 249308 534653 249317 534771
rect 175851 533590 175860 533730
rect 176000 533590 176009 533730
rect 101784 530884 101940 530889
rect 27853 530586 27862 530646
rect 27922 530630 27931 530646
rect 27922 530602 29220 530630
rect 27922 530586 27931 530602
rect 29350 530566 29378 530722
rect 102490 530568 102518 530990
rect 175860 530902 176000 533590
rect 175906 530560 175934 530902
rect 249190 530862 249308 534653
rect 322604 530890 322746 535759
rect 249230 530562 249258 530862
rect 322646 530560 322674 530890
rect 395928 530802 396042 536843
rect 542593 531406 542602 531466
rect 542662 531406 542671 531466
rect 469341 530970 469350 531060
rect 469440 530970 469449 531060
rect 395970 530562 395998 530802
rect 469350 530786 469440 530970
rect 469386 530564 469414 530786
rect 542618 530566 542646 531406
rect 552899 530658 552989 530667
rect 543074 530630 552899 530658
rect 542772 530602 552899 530630
rect 543074 530568 552899 530602
rect 552899 530559 552989 530568
rect 27649 500394 27658 500454
rect 27718 500438 27727 500454
rect 27718 500410 29214 500438
rect 27718 500394 27727 500410
rect 27649 470202 27658 470262
rect 27718 470246 27727 470262
rect 27718 470218 29214 470246
rect 27718 470202 27727 470218
rect 27649 440010 27658 440070
rect 27718 440054 27727 440070
rect 27718 440026 29214 440054
rect 27718 440010 27727 440026
rect 27649 409886 27658 409946
rect 27718 409930 27727 409946
rect 27718 409902 29214 409930
rect 27718 409886 27727 409902
rect 27649 379694 27658 379754
rect 27718 379738 27727 379754
rect 27718 379710 29214 379738
rect 27718 379694 27727 379710
rect 27649 349502 27658 349562
rect 27718 349546 27727 349562
rect 27718 349518 29214 349546
rect 27718 349502 27727 349518
rect 27649 319378 27658 319438
rect 27718 319422 27727 319438
rect 27718 319394 29214 319422
rect 27718 319378 27727 319394
rect 26112 295425 26699 295527
rect 26801 295425 27404 295527
rect 26112 295414 27404 295425
rect 26586 289246 26646 289255
rect 26646 289202 29214 289230
rect 26586 289177 26646 289186
rect 555728 274218 555788 274227
rect 542778 274174 555728 274202
rect 555728 274149 555788 274158
rect 26818 259054 26878 259063
rect 26878 259010 29212 259038
rect 26818 258985 26878 258994
rect 14310 248857 14603 248959
rect 14705 248857 14978 248959
rect 14310 248824 14978 248857
rect 27056 228862 27116 228871
rect 27116 228818 29220 228846
rect 27056 228793 27116 228802
rect 27284 198738 27344 198747
rect 27344 198694 29214 198722
rect 27284 198669 27344 198678
rect 27518 168546 27578 168555
rect 27578 168502 29212 168530
rect 27518 168477 27578 168486
rect 27752 138354 27812 138363
rect 27812 138310 29210 138338
rect 27752 138285 27812 138294
rect 9596 121235 9995 121337
rect 10097 121235 10498 121337
rect 9596 121187 10498 121235
rect 27976 108230 28036 108239
rect 28036 108186 29216 108214
rect 27976 108161 28036 108170
rect 6634 81559 7165 81661
rect 7267 81559 7768 81661
rect 6634 81555 7768 81559
rect 28230 78038 28290 78047
rect 28290 77994 29214 78022
rect 28230 77969 28290 77978
rect 567378 48203 567972 662985
rect 569844 662044 570372 662048
rect 569839 662039 580601 662044
rect 569839 661511 569844 662039
rect 570372 661511 580601 662039
rect 569839 661506 580601 661511
rect 569844 661502 570372 661506
rect 580063 92861 580601 661506
rect 580063 92759 580277 92861
rect 580379 92759 580601 92861
rect 580063 92707 580601 92759
rect 567378 48101 567603 48203
rect 567705 48101 567972 48203
rect 567378 48091 567972 48101
rect 28522 47846 28582 47855
rect 28582 47802 29220 47830
rect 28522 47777 28582 47786
rect 28864 17722 28924 17731
rect 558978 17722 559038 17731
rect 28924 17678 29230 17706
rect 542780 17678 558978 17706
rect 28864 17653 28924 17662
rect 558978 17653 559038 17662
rect 579052 14662 579174 14668
rect 578190 14540 578199 14662
rect 578321 14540 579052 14662
rect 578575 9936 578697 14540
rect 579052 14534 579174 14540
rect 580143 14662 580265 14668
rect 582049 14658 582151 14662
rect 580265 14653 582156 14658
rect 580265 14551 582049 14653
rect 582151 14551 582156 14653
rect 580265 14546 582156 14551
rect 582049 14542 582151 14546
rect 580143 14534 580265 14540
rect 579064 9936 579186 9942
rect 578575 9814 579064 9936
rect 578575 5206 578697 9814
rect 579064 9808 579186 9814
rect 580155 9936 580277 9942
rect 582061 9932 582163 9936
rect 580277 9927 582168 9932
rect 580277 9825 582061 9927
rect 582163 9825 582168 9927
rect 580277 9820 582168 9825
rect 582061 9816 582163 9820
rect 580155 9808 580277 9814
rect 579176 5206 579298 5212
rect 578575 5084 579176 5206
rect 578575 5075 578697 5084
rect 579176 5078 579298 5084
rect 580267 5206 580389 5212
rect 582173 5202 582275 5206
rect 580389 5197 582280 5202
rect 580389 5095 582173 5197
rect 582275 5095 582280 5197
rect 580389 5090 582280 5095
rect 582173 5086 582275 5090
rect 580267 5078 580389 5084
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 171904 701992 172024 702112
rect 174410 701992 174530 702112
rect 223692 701992 223812 702112
rect 226092 701992 226212 702112
rect 325330 701992 325450 702112
rect 327840 701992 327960 702112
rect 26120 700222 26580 700682
rect 18310 697260 18730 697680
rect 28697 697220 29117 697640
rect 30193 694278 30603 694688
rect 9732 685550 10132 685950
rect 2919 682546 3223 682850
rect 9010 679566 9410 679966
rect 133170 698890 133538 699258
rect 122377 698407 122827 698857
rect 130731 698423 131181 698873
rect 70569 697301 70947 697679
rect 78989 697275 79367 697653
rect 81985 695439 82391 695845
rect 122466 695406 122834 695774
rect 71597 694264 72003 694670
rect 69181 690163 69599 690581
rect 171904 699020 172024 699140
rect 196540 700255 197122 700837
rect 174410 699030 174514 699134
rect 194112 697430 194572 697890
rect 186408 695068 186788 695448
rect 185244 694488 185388 694632
rect 134489 690165 134915 690591
rect 12317 679561 12727 679971
rect 4127 656495 5109 657477
rect 9596 658559 10498 659461
rect 7866 549131 8170 549435
rect 11763 654311 12653 655201
rect 9895 600461 10093 600659
rect 4603 338647 4705 338749
rect 7079 548373 7421 548715
rect 9963 547309 10213 547559
rect 90758 622092 90818 622152
rect 90674 619916 90734 619976
rect 90962 617672 91022 617732
rect 90760 615428 90820 615488
rect 90750 613184 90810 613244
rect 90708 611008 90768 611068
rect 90732 608764 90792 608824
rect 90666 606520 90726 606580
rect 90700 604276 90760 604336
rect 12237 381869 12339 381971
rect 14575 601153 14781 601359
rect 14573 550011 14823 550261
rect 16898 596625 17238 596965
rect 74702 601222 74762 601282
rect 98678 619880 98798 620000
rect 98365 617659 98483 617777
rect 98061 615403 98179 615521
rect 97757 613145 97875 613263
rect 97467 610937 97585 611055
rect 97187 608739 97305 608857
rect 96883 606483 97001 606601
rect 82522 600526 82582 600586
rect 74050 594444 74167 594561
rect 91824 596740 91936 596852
rect 96629 604249 96747 604367
rect 96634 594150 96742 594258
rect 96888 593854 96996 593962
rect 97192 593586 97300 593694
rect 97472 593316 97580 593424
rect 97762 593004 97870 593112
rect 98066 592714 98174 592822
rect 98370 592424 98478 592532
rect 185658 693166 185794 693302
rect 185271 617597 185361 617687
rect 219627 699849 220101 700323
rect 210649 695073 211019 695443
rect 221404 698892 221768 699256
rect 223696 699044 223800 699148
rect 264688 700300 264872 700484
rect 226094 699064 226198 699168
rect 209714 693586 210102 693974
rect 204962 692052 205298 692388
rect 202461 686458 202807 686804
rect 313069 700141 313737 700809
rect 321259 700150 321924 700815
rect 310807 698891 311169 699253
rect 314732 697572 315200 698040
rect 325346 699004 325450 699108
rect 327840 699016 327944 699120
rect 323712 696231 324526 697045
rect 282157 663213 282311 663367
rect 279759 661640 279819 661700
rect 215183 656787 215421 657025
rect 215886 654524 216138 654776
rect 222630 648298 222758 648426
rect 220299 638769 220389 638859
rect 220155 634239 220245 634329
rect 294492 640050 294552 640110
rect 285236 633906 285428 634098
rect 267177 632565 267379 632767
rect 244672 628506 244856 628690
rect 265750 628502 265934 628686
rect 245670 628155 245872 628357
rect 285231 632277 285433 632479
rect 282616 631830 282716 631930
rect 289037 631835 289127 631925
rect 294053 629755 294299 630001
rect 291980 629376 292080 629476
rect 267182 628160 267374 628352
rect 291985 626745 292075 626835
rect 294822 626519 295332 627029
rect 245715 625651 245805 625741
rect 294048 625504 294304 625760
rect 292225 623651 292315 623741
rect 294316 623646 294416 623746
rect 185681 617583 185771 617673
rect 186413 617369 186783 617739
rect 182728 615814 182828 615914
rect 183066 615408 183166 615508
rect 183071 607593 183161 607683
rect 182733 605609 182823 605699
rect 270579 595293 270669 595383
rect 98683 592153 98793 592263
rect 90325 585619 90415 585709
rect 90322 578311 90427 578416
rect 90690 568566 90750 568626
rect 90978 566322 91038 566382
rect 90776 564078 90836 564138
rect 90766 561834 90826 561894
rect 90724 559658 90784 559718
rect 90748 557414 90808 557474
rect 90682 555170 90742 555230
rect 90716 552926 90776 552986
rect 93700 578306 93815 578421
rect 17053 468313 17155 468415
rect 22543 543995 22797 544249
rect 29318 541694 29423 541799
rect 22621 425091 22723 425193
rect 26511 539055 26957 539501
rect 29312 534202 29416 534306
rect 74718 550110 74778 550170
rect 82538 547410 82598 547470
rect 91840 544072 91952 544184
rect 90331 541689 90446 541804
rect 101784 567946 101940 568102
rect 101363 566283 101521 566441
rect 100896 564030 101060 564194
rect 100463 561799 100593 561929
rect 99970 559604 100090 559724
rect 99470 557376 99598 557504
rect 99053 555135 99187 555269
rect 98621 552889 98755 553023
rect 93705 541694 93810 541799
rect 74319 533069 74430 533180
rect 98626 532810 98750 532934
rect 99058 532560 99182 532684
rect 99475 532319 99593 532437
rect 99975 532105 100085 532215
rect 100468 531840 100588 531960
rect 100901 531531 101055 531685
rect 101368 531202 101516 531350
rect 183933 561543 184023 561633
rect 149945 556583 150035 556673
rect 149545 554599 149635 554689
rect 149540 549262 149640 549362
rect 251836 557474 251896 557534
rect 226891 555063 227077 555249
rect 182912 550926 183012 551026
rect 149940 548518 150040 548618
rect 226886 552270 227082 552466
rect 326104 692323 327354 693573
rect 323930 550819 324238 551127
rect 417389 698907 417731 699249
rect 403319 696236 404123 697040
rect 414474 696236 415278 697040
rect 470545 698901 470899 699255
rect 459850 695870 460194 696214
rect 456956 692760 457524 693328
rect 467602 692760 468170 693328
rect 401679 690713 402065 691099
rect 562836 695304 563216 695684
rect 562085 692161 562779 692855
rect 569177 692179 569871 692873
rect 560028 689348 560392 689712
rect 333298 683126 334002 683830
rect 572986 680148 573554 680716
rect 580556 680148 581124 680716
rect 567394 662985 567978 663569
rect 545439 632909 546229 633699
rect 333303 631453 333997 632147
rect 332404 626524 332904 627024
rect 330329 625231 331051 625953
rect 330324 617290 331056 618022
rect 332399 612509 332909 613019
rect 545434 582000 546234 582800
rect 225796 548492 225916 548612
rect 326375 548281 326869 548775
rect 102444 547371 102574 547501
rect 101789 530889 101935 531035
rect 395928 536843 396042 536957
rect 322604 535759 322746 535901
rect 249190 534653 249308 534771
rect 175860 533590 176000 533730
rect 27862 530586 27922 530646
rect 542602 531406 542662 531466
rect 469350 530970 469440 531060
rect 552899 530568 552989 530658
rect 27658 500394 27718 500454
rect 27658 470202 27718 470262
rect 27658 440010 27718 440070
rect 27658 409886 27718 409946
rect 27658 379694 27718 379754
rect 27658 349502 27718 349562
rect 27658 319378 27718 319438
rect 26699 295425 26801 295527
rect 26586 289186 26646 289246
rect 555728 274158 555788 274218
rect 26818 258994 26878 259054
rect 14603 248857 14705 248959
rect 27056 228802 27116 228862
rect 27284 198678 27344 198738
rect 27518 168486 27578 168546
rect 27752 138294 27812 138354
rect 9995 121235 10097 121337
rect 27976 108170 28036 108230
rect 7165 81559 7267 81661
rect 28230 77978 28290 78038
rect 569844 661511 570372 662039
rect 580277 92759 580379 92861
rect 567603 48101 567705 48203
rect 28522 47786 28582 47846
rect 28864 17662 28924 17722
rect 558978 17662 559038 17722
rect 578199 14540 578321 14662
rect 582049 14551 582151 14653
rect 582061 9825 582163 9927
rect 582173 5095 582275 5197
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 18305 697680 18735 702300
rect 26115 700682 26585 700687
rect 26115 700222 26120 700682
rect 26580 700222 26585 700682
rect 26115 700217 26585 700222
rect 18305 697260 18310 697680
rect 18730 697260 18735 697680
rect 18305 697255 18735 697260
rect 26120 691015 26580 700217
rect 70564 697679 70952 702300
rect 122372 698857 122832 702300
rect 167845 700837 168427 702300
rect 171820 702112 172132 702300
rect 171820 701992 171904 702112
rect 172024 701992 172132 702112
rect 171820 701948 172132 701992
rect 174326 702112 174638 702300
rect 174326 701992 174410 702112
rect 174530 701992 174638 702112
rect 174326 701948 174638 701992
rect 178141 700837 178723 702300
rect 196535 700837 197127 700842
rect 167845 700255 196540 700837
rect 197122 700255 197127 700837
rect 219622 700340 220106 702300
rect 223608 702112 223920 702300
rect 223608 701992 223692 702112
rect 223812 701992 223920 702112
rect 223608 701948 223920 701992
rect 226008 702112 226320 702300
rect 226008 701992 226092 702112
rect 226212 701992 226320 702112
rect 226008 701948 226320 701992
rect 229792 700340 230276 702300
rect 321251 701312 321929 702300
rect 325246 702112 325558 702300
rect 325246 701992 325330 702112
rect 325450 701992 325558 702112
rect 325246 701948 325558 701992
rect 327756 702112 328068 702300
rect 327756 701992 327840 702112
rect 327960 701992 328068 702112
rect 327756 701948 328068 701992
rect 321254 700815 321929 701312
rect 196535 700250 197127 700255
rect 219588 700323 230276 700340
rect 219588 699872 219627 700323
rect 219622 699849 219627 699872
rect 220101 699872 230276 700323
rect 264508 700809 313742 700814
rect 264508 700484 313069 700809
rect 264508 700300 264688 700484
rect 264872 700300 313069 700484
rect 264508 700141 313069 700300
rect 313737 700141 313742 700809
rect 264508 700136 313742 700141
rect 321254 700150 321259 700815
rect 321924 700814 321929 700815
rect 331423 700814 332101 702300
rect 321924 700150 332101 700814
rect 321254 700136 332101 700150
rect 220101 699849 220106 699872
rect 220606 699856 230276 699872
rect 219622 699844 220106 699849
rect 132958 699258 412641 699376
rect 132958 698890 133170 699258
rect 133538 699256 412641 699258
rect 133538 699140 221404 699256
rect 133538 699020 171904 699140
rect 172024 699134 221404 699140
rect 172024 699030 174410 699134
rect 174514 699030 221404 699134
rect 172024 699020 221404 699030
rect 133538 698892 221404 699020
rect 221768 699253 412641 699256
rect 221768 699168 310807 699253
rect 221768 699148 226094 699168
rect 221768 699044 223696 699148
rect 223800 699064 226094 699148
rect 226198 699064 310807 699168
rect 223800 699044 310807 699064
rect 221768 698892 310807 699044
rect 133538 698891 310807 698892
rect 311169 699120 412641 699253
rect 311169 699108 327840 699120
rect 311169 699004 325346 699108
rect 325450 699016 327840 699108
rect 327944 699016 412641 699120
rect 325450 699004 412641 699016
rect 311169 698891 412641 699004
rect 133538 698890 412641 698891
rect 122372 698407 122377 698857
rect 122827 698407 122832 698857
rect 122372 698402 122832 698407
rect 130726 698873 131186 698878
rect 130726 698423 130731 698873
rect 131181 698423 131186 698873
rect 132958 698770 412641 698890
rect 413247 698770 413253 699376
rect 28692 697640 29122 697665
rect 28692 697220 28697 697640
rect 29117 697220 29122 697640
rect 70564 697301 70569 697679
rect 70947 697301 70952 697679
rect 130726 697890 131186 698423
rect 314727 698040 315205 698045
rect 194107 697890 194577 697895
rect 70564 697296 70952 697301
rect 78984 697653 79372 697658
rect 28692 693414 29122 697220
rect 78984 697275 78989 697653
rect 79367 697275 79372 697653
rect 130726 697430 194112 697890
rect 194572 697430 194577 697890
rect 314727 697572 314732 698040
rect 315200 697572 315205 698040
rect 314727 697567 315205 697572
rect 194107 697425 194577 697430
rect 30008 694688 72188 694840
rect 30008 694278 30193 694688
rect 30603 694670 72188 694688
rect 30603 694278 71597 694670
rect 30008 694264 71597 694278
rect 72003 694264 72188 694670
rect 78984 694756 79372 697275
rect 81812 695845 122960 696102
rect 81812 695439 81985 695845
rect 82391 695774 122960 695845
rect 82391 695439 122466 695774
rect 81812 695406 122466 695439
rect 122834 695406 122960 695774
rect 81812 695194 122960 695406
rect 186403 695448 186793 695453
rect 186403 695068 186408 695448
rect 186788 695443 211024 695448
rect 186788 695073 210649 695443
rect 211019 695073 211024 695443
rect 186788 695068 211024 695073
rect 186403 695063 186793 695068
rect 78984 694632 185462 694756
rect 78984 694488 185244 694632
rect 185388 694488 185462 694632
rect 78984 694368 185462 694488
rect 30008 693984 72188 694264
rect 209709 693974 210107 693979
rect 209709 693586 209714 693974
rect 210102 693586 210107 693974
rect 209709 693581 210107 693586
rect 28692 693302 185918 693414
rect 28692 693166 185658 693302
rect 185794 693166 185918 693302
rect 28692 692984 185918 693166
rect 204957 692388 205303 692393
rect 204957 692052 204962 692388
rect 205298 692052 205303 692388
rect 67914 691015 183014 691032
rect 15173 690814 183014 691015
rect 15173 689916 30406 690814
rect 34854 690591 183014 690814
rect 34854 690581 134489 690591
rect 34854 690163 69181 690581
rect 69599 690165 134489 690581
rect 134915 690165 183014 690591
rect 69599 690163 183014 690165
rect 34854 689916 183014 690163
rect 15173 689748 183014 689916
rect 9727 685950 10137 685955
rect 15173 685950 16440 689748
rect 67914 689708 183014 689748
rect 9727 685550 9732 685950
rect 10132 685550 16466 685950
rect 9727 685545 10137 685550
rect -800 682855 1700 685242
rect 181690 683002 183014 689708
rect 202456 686804 202812 686809
rect 204957 686804 205303 692052
rect 209714 687274 210102 693581
rect 314732 687274 315200 697567
rect 323707 697045 324531 697050
rect 415421 697045 416235 702300
rect 417384 699254 417736 699260
rect 417384 698907 417389 698912
rect 417731 698907 417736 698912
rect 417384 698902 417736 698907
rect 323707 696231 323712 697045
rect 324526 697040 404128 697045
rect 324526 696236 403319 697040
rect 404123 696236 404128 697040
rect 324526 696231 404128 696236
rect 414450 697040 416235 697045
rect 414450 696236 414474 697040
rect 415278 696236 416235 697040
rect 414450 696231 416235 696236
rect 323707 696226 324531 696231
rect 459845 696214 460199 696219
rect 459845 695870 459850 696214
rect 460194 695870 460199 696214
rect 459845 695865 460199 695870
rect 326099 693573 327359 693578
rect 326099 692323 326104 693573
rect 327354 693328 457696 693573
rect 327354 692760 456956 693328
rect 457524 692760 457696 693328
rect 327354 692323 457696 692760
rect 326099 692318 327359 692323
rect 401674 691099 402070 691104
rect 401674 690713 401679 691099
rect 402065 690713 402070 691099
rect 401674 690708 402070 690713
rect 401679 687274 402065 690708
rect 459850 687274 460194 695865
rect 467273 693328 468523 702300
rect 470540 699260 470904 699266
rect 470540 698901 470545 698906
rect 470899 698901 470904 698906
rect 470540 698896 470904 698901
rect 512816 699204 515276 702340
rect 520594 699204 523054 702340
rect 566594 702300 571594 704800
rect 467273 692760 467602 693328
rect 468170 692760 468523 693328
rect 467273 692705 468523 692760
rect 512816 696744 520568 699204
rect 523028 696744 523054 699204
rect 512816 695086 515276 696744
rect 512816 692620 515276 692626
rect 555818 695684 563468 696048
rect 555818 695304 562836 695684
rect 563216 695304 563468 695684
rect 555818 694724 563468 695304
rect 555818 687274 557142 694724
rect 569172 692873 569876 702300
rect 562080 692855 562784 692860
rect 562080 692161 562085 692855
rect 562779 692161 562784 692855
rect 569172 692179 569177 692873
rect 569871 692179 569876 692873
rect 569172 692174 569876 692179
rect 560023 689717 560397 689723
rect 560023 689348 560028 689353
rect 560392 689348 560397 689353
rect 560023 689343 560397 689348
rect 202456 686458 202461 686804
rect 202807 686458 205303 686804
rect 202456 686453 202812 686458
rect 207618 685950 557142 687274
rect 207618 683002 208942 685950
rect 333293 683830 334007 683835
rect 562080 683830 562784 692161
rect 333293 683126 333298 683830
rect 334002 683126 562784 683830
rect 333293 683121 334007 683126
rect -800 682850 3228 682855
rect -800 682546 2919 682850
rect 3223 682546 3228 682850
rect -800 682541 3228 682546
rect -800 680242 1700 682541
rect 181690 681678 208942 683002
rect 582300 680761 584800 682984
rect 572285 680716 573670 680761
rect 572285 680148 572986 680716
rect 573554 680148 573670 680716
rect 572285 680039 573670 680148
rect 580494 680716 584800 680761
rect 580494 680148 580556 680716
rect 581124 680148 584800 680716
rect 580494 680039 584800 680148
rect 12312 679971 12732 679976
rect 9005 679966 12317 679971
rect 9005 679566 9010 679966
rect 9410 679566 12317 679966
rect 9005 679561 12317 679566
rect 12727 679561 12732 679971
rect 12312 679556 12732 679561
rect 282128 663569 567983 663574
rect 282128 663367 567394 663569
rect 282128 663213 282157 663367
rect 282311 663213 567394 663367
rect 282128 662985 567394 663213
rect 567978 662985 567983 663569
rect 282128 662980 567983 662985
rect 279734 662039 570377 662044
rect 279734 661700 569844 662039
rect 279734 661640 279759 661700
rect 279819 661640 569844 661700
rect 279734 661511 569844 661640
rect 570372 661511 570377 662039
rect 279734 661506 570377 661511
rect 9475 659461 222804 659540
rect 9475 658559 9596 659461
rect 10498 658559 222804 659461
rect 9475 658398 222804 658559
rect 4122 657477 215506 657482
rect 4122 656495 4127 657477
rect 5109 657025 215506 657477
rect 5109 656787 215183 657025
rect 215421 656787 215506 657025
rect 5109 656495 215506 656787
rect 4122 656490 215506 656495
rect 11758 655201 216158 655206
rect 11758 654311 11763 655201
rect 12653 654776 216158 655201
rect 12653 654524 215886 654776
rect 216138 654524 216158 654776
rect 12653 654311 216158 654524
rect 11758 654306 216158 654311
rect -800 648564 1660 648642
rect -800 643900 15002 648564
rect 19666 643900 19672 648564
rect 222572 648426 222802 658398
rect 222572 648298 222630 648426
rect 222758 648298 222802 648426
rect 222572 648260 222802 648298
rect -800 643842 1660 643900
rect -800 638558 1660 638642
rect 8408 638558 13072 643900
rect 294472 640110 297043 640136
rect 294472 640050 294492 640110
rect 294552 640050 297043 640110
rect 294472 639998 297043 640050
rect 220294 638859 220600 638864
rect 220294 638769 220299 638859
rect 220389 638769 220600 638859
rect 220294 638764 220600 638769
rect -800 633894 13072 638558
rect 220150 634329 220420 634334
rect 220150 634239 220155 634329
rect 220245 634239 220420 634329
rect 220150 634234 220420 634239
rect 281465 634098 285433 634103
rect 281465 633906 285236 634098
rect 285428 633906 285433 634098
rect 281465 633901 285433 633906
rect -800 633842 1660 633894
rect 267172 632767 267384 632772
rect 281465 632767 281667 633901
rect 296905 633393 297043 639998
rect 321650 633699 546234 633704
rect 321650 633393 545439 633699
rect 296905 633255 545439 633393
rect 321650 632909 545439 633255
rect 546229 632909 546234 633699
rect 321650 632904 546234 632909
rect 267172 632565 267177 632767
rect 267379 632565 281667 632767
rect 267172 632560 267384 632565
rect 285226 632479 285438 632484
rect 285226 632277 285231 632479
rect 285433 632277 289887 632479
rect 285226 632272 285438 632277
rect 282611 631930 282721 631935
rect 282611 631830 282616 631930
rect 282716 631925 289132 631930
rect 282716 631835 289037 631925
rect 289127 631835 289132 631925
rect 282716 631830 289132 631835
rect 289685 631921 289887 632277
rect 329060 632147 334076 632152
rect 329060 631921 333303 632147
rect 282611 631825 282721 631830
rect 289685 631719 333303 631921
rect 270312 631406 289469 631592
rect 329060 631453 333303 631719
rect 333997 631453 334076 632147
rect 329060 631448 334076 631453
rect 270314 628860 270414 631406
rect 289283 630453 289469 631406
rect 572285 630692 573007 680039
rect 582300 677984 584800 680039
rect 582340 644550 584800 644584
rect 575932 639830 575938 644550
rect 580658 639830 584800 644550
rect 328964 630453 573007 630692
rect 577382 632996 579842 639830
rect 582340 639784 584800 639830
rect 582340 632996 584800 634584
rect 577382 630536 584800 632996
rect 289283 630267 573007 630453
rect 292322 630001 294304 630006
rect 292322 629928 294053 630001
rect 288724 629828 294053 629928
rect 292322 629755 294053 629828
rect 294299 629755 294304 630001
rect 328964 629970 573007 630267
rect 582340 629784 584800 630536
rect 292322 629750 294304 629755
rect 291952 629476 328227 629556
rect 291952 629376 291980 629476
rect 292080 629376 328227 629476
rect 291952 629310 328227 629376
rect 244667 628690 244861 628695
rect 265745 628690 265939 628691
rect 244667 628506 244672 628690
rect 244856 628686 265950 628690
rect 244856 628506 265750 628686
rect 244667 628501 244861 628506
rect 265745 628502 265750 628506
rect 265934 628506 265950 628686
rect 265934 628502 265939 628506
rect 265745 628497 265939 628502
rect 327981 628382 328227 629310
rect 245665 628357 245877 628362
rect 245665 628155 245670 628357
rect 245872 628352 267379 628357
rect 245872 628160 267182 628352
rect 267374 628160 267379 628352
rect 245872 628155 267379 628160
rect 245665 628150 245877 628155
rect 327981 627637 577818 628382
rect 328008 627634 577818 627637
rect 294817 627029 295337 627034
rect 268576 626835 292080 626840
rect 268576 626745 291985 626835
rect 292075 626745 292080 626835
rect 268576 626740 292080 626745
rect 294817 626519 294822 627029
rect 295332 627024 332909 627029
rect 295332 626524 332404 627024
rect 332904 626524 332909 627024
rect 295332 626519 332909 626524
rect 294817 626514 295337 626519
rect 294006 625953 331056 625958
rect 294006 625760 330329 625953
rect 245710 625741 245810 625746
rect 245710 625651 245715 625741
rect 245805 625651 245810 625741
rect 245710 625646 245810 625651
rect 294006 625504 294048 625760
rect 294304 625504 330329 625760
rect 294006 625231 330329 625504
rect 331051 625231 331056 625953
rect 294006 625226 331056 625231
rect 294290 623746 574212 623952
rect 292048 623741 292320 623746
rect 292048 623651 292225 623741
rect 292315 623651 292320 623741
rect 292048 623646 292320 623651
rect 294290 623646 294316 623746
rect 294416 623646 574212 623746
rect 294290 623396 574212 623646
rect 90730 622152 93205 622204
rect 90730 622092 90758 622152
rect 90818 622092 93205 622152
rect 90730 622054 93205 622092
rect 93055 620431 93205 622054
rect 292480 621874 292580 623004
rect 292476 621228 569437 621874
rect 93055 620281 137841 620431
rect 137991 620281 137997 620431
rect 140292 620430 140440 620436
rect 140292 620276 140440 620282
rect 90649 620000 137091 620037
rect 90649 619976 98678 620000
rect 90649 619916 90674 619976
rect 90734 619916 98678 619976
rect 90649 619880 98678 619916
rect 98798 619880 137091 620000
rect 90649 619859 137091 619880
rect 90925 617777 135727 617803
rect 90925 617732 98365 617777
rect 90925 617672 90962 617732
rect 91022 617672 98365 617732
rect 90925 617659 98365 617672
rect 98483 617659 135727 617777
rect 90925 617625 135727 617659
rect 90737 615521 134349 615543
rect 90737 615488 98061 615521
rect 90737 615428 90760 615488
rect 90820 615428 98061 615488
rect 90737 615403 98061 615428
rect 98179 615403 134349 615521
rect 90737 615365 134349 615403
rect 90723 613263 132889 613299
rect 90723 613244 97757 613263
rect 90723 613184 90750 613244
rect 90810 613184 97757 613244
rect 90723 613145 97757 613184
rect 97875 613145 132889 613263
rect 90723 613121 132889 613145
rect 90679 611068 131559 611103
rect 90679 611008 90708 611068
rect 90768 611055 131559 611068
rect 90768 611008 97467 611055
rect 90679 610937 97467 611008
rect 97585 610937 131559 611055
rect 90679 610925 131559 610937
rect 90707 608857 130513 608885
rect 90707 608824 97187 608857
rect 90707 608764 90732 608824
rect 90792 608764 97187 608824
rect 90707 608739 97187 608764
rect 97305 608739 130513 608857
rect 90707 608707 130513 608739
rect 90647 606601 129595 606637
rect 90647 606600 96883 606601
rect 90646 606580 96883 606600
rect 90646 606520 90666 606580
rect 90726 606520 96883 606580
rect 90646 606504 96883 606520
rect 90647 606483 96883 606504
rect 97001 606483 129595 606601
rect 90647 606459 129595 606483
rect 90677 604367 128845 604395
rect 90677 604336 96629 604367
rect 90677 604276 90700 604336
rect 90760 604276 96629 604336
rect 90677 604249 96629 604276
rect 96747 604249 128845 604367
rect 90677 604217 128845 604249
rect 128667 602614 128845 604217
rect 129417 602912 129595 606459
rect 130335 603190 130513 608707
rect 131381 603472 131559 610925
rect 132711 603774 132889 613121
rect 134171 604048 134349 615365
rect 135549 604364 135727 617625
rect 136913 604652 137091 619859
rect 330319 618022 331061 618027
rect 186408 617739 186788 617744
rect 185266 617687 185366 617692
rect 185266 617597 185271 617687
rect 185361 617597 185366 617687
rect 182723 615914 182833 615919
rect 185266 615914 185366 617597
rect 182723 615814 182728 615914
rect 182828 615814 185366 615914
rect 185676 617673 185776 617678
rect 185676 617583 185681 617673
rect 185771 617583 185776 617673
rect 182723 615809 182833 615814
rect 183061 615508 183171 615513
rect 185676 615508 185776 617583
rect 183061 615408 183066 615508
rect 183166 615408 185776 615508
rect 186408 617369 186413 617739
rect 186783 617369 186788 617739
rect 183061 615403 183171 615408
rect 186408 612782 186788 617369
rect 330319 617290 330324 618022
rect 331056 617290 563858 618022
rect 330319 617285 331061 617290
rect 181778 612402 186788 612782
rect 332352 613019 558426 613476
rect 332352 612509 332399 613019
rect 332909 612509 558426 613019
rect 332352 611640 558426 612509
rect 181472 607683 183166 607688
rect 181472 607593 183071 607683
rect 183161 607593 183166 607683
rect 181472 607588 183166 607593
rect 181192 605699 182828 605704
rect 181192 605609 182733 605699
rect 182823 605609 182828 605699
rect 181192 605604 182828 605609
rect 136913 604474 142902 604652
rect 135549 604186 142904 604364
rect 134171 603870 142912 604048
rect 132711 603596 142914 603774
rect 131381 603294 142898 603472
rect 130335 603012 142894 603190
rect 129417 602734 142912 602912
rect 128667 602436 142914 602614
rect 14570 601359 74802 601364
rect 14570 601153 14575 601359
rect 14781 601282 74802 601359
rect 14781 601222 74702 601282
rect 74762 601222 74802 601282
rect 14781 601153 74802 601222
rect 14570 601148 74802 601153
rect 9890 600659 82612 600664
rect 9890 600461 9895 600659
rect 10093 600586 82612 600659
rect 10093 600526 82522 600586
rect 82582 600526 82612 600586
rect 10093 600461 82612 600526
rect 9890 600456 82612 600461
rect 16893 596965 91972 596970
rect 16893 596625 16898 596965
rect 17238 596852 91972 596965
rect 17238 596740 91824 596852
rect 91936 596740 91972 596852
rect 17238 596625 91972 596740
rect 16893 596620 91972 596625
rect 270283 595383 270674 595388
rect 270283 595293 270579 595383
rect 270669 595293 270674 595383
rect 270283 595288 270674 595293
rect 24254 594565 24386 594570
rect 74045 594565 74172 594566
rect 24253 594564 74179 594565
rect 24253 594432 24254 594564
rect 24386 594561 74179 594564
rect 24386 594444 74050 594561
rect 74167 594444 74179 594561
rect 24386 594432 74179 594444
rect 24253 594431 74179 594432
rect 24254 594426 24386 594431
rect 24594 594263 24710 594268
rect 24593 594262 96747 594263
rect 24593 594146 24594 594262
rect 24710 594258 96747 594262
rect 24710 594150 96634 594258
rect 96742 594150 96747 594258
rect 24710 594146 96747 594150
rect 24593 594145 96747 594146
rect 24594 594140 24710 594145
rect 24914 593967 25030 593972
rect 24913 593966 97001 593967
rect 24913 593850 24914 593966
rect 25030 593962 97001 593966
rect 25030 593854 96888 593962
rect 96996 593854 97001 593962
rect 25030 593850 97001 593854
rect 24913 593849 97001 593850
rect 24914 593844 25030 593849
rect 25216 593699 25332 593704
rect 25215 593698 97305 593699
rect 25215 593582 25216 593698
rect 25332 593694 97305 593698
rect 25332 593586 97192 593694
rect 97300 593586 97305 593694
rect 25332 593582 97305 593586
rect 25215 593581 97305 593582
rect 25216 593576 25332 593581
rect 25494 593429 25610 593434
rect 25493 593428 97585 593429
rect 25493 593312 25494 593428
rect 25610 593424 97585 593428
rect 25610 593316 97472 593424
rect 97580 593316 97585 593424
rect 25610 593312 97585 593316
rect 25493 593311 97585 593312
rect 25494 593306 25610 593311
rect 25784 593117 25900 593122
rect 25783 593116 97875 593117
rect 25783 593000 25784 593116
rect 25900 593112 97875 593116
rect 25900 593004 97762 593112
rect 97870 593004 97875 593112
rect 25900 593000 97875 593004
rect 25783 592999 97875 593000
rect 25784 592994 25900 592999
rect 26066 592827 26182 592832
rect 26065 592826 98179 592827
rect 26065 592710 26066 592826
rect 26182 592822 98179 592826
rect 26182 592714 98066 592822
rect 98174 592714 98179 592822
rect 26182 592710 98179 592714
rect 26065 592709 98179 592710
rect 26066 592704 26182 592709
rect 26318 592537 26434 592542
rect 26317 592536 98483 592537
rect 26317 592420 26318 592536
rect 26434 592532 98483 592536
rect 26434 592424 98370 592532
rect 98478 592424 98483 592532
rect 26434 592420 98483 592424
rect 26317 592419 98483 592420
rect 26318 592414 26434 592419
rect 26555 592268 26673 592273
rect 26554 592267 98798 592268
rect 26554 592149 26555 592267
rect 26673 592263 98798 592267
rect 26673 592153 98683 592263
rect 98793 592153 98798 592263
rect 26673 592149 98798 592153
rect 26554 592148 98798 592149
rect 26555 592143 26673 592148
rect 270283 588060 270478 595288
rect 270282 588052 548702 588060
rect 270282 587608 552174 588052
rect 90320 585709 94722 585714
rect 90320 585619 90325 585709
rect 90415 585619 94722 585709
rect 90320 585614 94722 585619
rect 544900 582800 547088 582992
rect 544900 582000 545434 582800
rect 546234 582000 547088 582800
rect 93695 578421 93820 578426
rect 90317 578416 93700 578421
rect 90317 578311 90322 578416
rect 90427 578311 93700 578416
rect 90317 578306 93700 578311
rect 93815 578306 93820 578421
rect 93695 578301 93820 578306
rect 90651 568626 90928 568687
rect 90651 568566 90690 568626
rect 90750 568566 90928 568626
rect 90651 568509 90928 568566
rect 90750 568121 90928 568509
rect 90750 568102 137107 568121
rect 90750 567946 101784 568102
rect 101940 567946 137107 568102
rect 90750 567943 137107 567946
rect 101779 567941 101945 567943
rect 90941 566441 135743 566453
rect 90941 566382 101363 566441
rect 90941 566322 90978 566382
rect 91038 566322 101363 566382
rect 90941 566283 101363 566322
rect 101521 566283 135743 566441
rect 90941 566275 135743 566283
rect -800 559442 1660 564242
rect 100891 564194 101065 564199
rect 100891 564193 100896 564194
rect 90753 564138 100896 564193
rect 90753 564078 90776 564138
rect 90836 564078 100896 564138
rect 90753 564030 100896 564078
rect 101060 564193 101065 564194
rect 101060 564030 134365 564193
rect 90753 564015 134365 564030
rect 90739 561929 132905 561949
rect 90739 561894 100463 561929
rect 90739 561834 90766 561894
rect 90826 561834 100463 561894
rect 90739 561799 100463 561834
rect 100593 561799 132905 561929
rect 90739 561771 132905 561799
rect 90695 559724 131575 559753
rect 90695 559718 99970 559724
rect 90695 559658 90724 559718
rect 90784 559658 99970 559718
rect 90695 559604 99970 559658
rect 100090 559604 131575 559724
rect 90695 559575 131575 559604
rect 90723 557525 99459 557535
rect 99742 557525 130529 557535
rect 90723 557504 130529 557525
rect 90723 557474 99470 557504
rect 90723 557414 90748 557474
rect 90808 557414 99470 557474
rect 90723 557376 99470 557414
rect 99598 557376 130529 557504
rect 90723 557366 130529 557376
rect 90723 557357 99459 557366
rect 99742 557357 130529 557366
rect 90663 555269 129611 555287
rect 90663 555250 99053 555269
rect 90662 555230 99053 555250
rect 90662 555170 90682 555230
rect 90742 555170 99053 555230
rect 90662 555154 99053 555170
rect 90663 555135 99053 555154
rect 99187 555135 129611 555269
rect 90663 555109 129611 555135
rect -800 549442 1660 554242
rect 90693 553023 128861 553045
rect 90693 552986 98621 553023
rect 90693 552926 90716 552986
rect 90776 552926 98621 552986
rect 90693 552889 98621 552926
rect 98755 552889 128861 553023
rect 90693 552867 128861 552889
rect 128683 551264 128861 552867
rect 129433 551562 129611 555109
rect 130351 551840 130529 557357
rect 131397 552122 131575 559575
rect 132727 552424 132905 561771
rect 134187 552698 134365 564015
rect 135565 553014 135743 566275
rect 136929 553302 137107 567943
rect 183928 561633 184028 561832
rect 183928 561543 183933 561633
rect 184023 561543 184028 561633
rect 183928 561538 184028 561543
rect 251770 557534 251966 557566
rect 251770 557474 251836 557534
rect 251896 557474 251966 557534
rect 149940 556673 150040 556678
rect 149940 556583 149945 556673
rect 150035 556583 150040 556673
rect 149940 556578 150040 556583
rect 226886 555852 250874 556048
rect 226886 555249 227082 555852
rect 250678 555744 250874 555852
rect 251770 555744 251966 557474
rect 250678 555548 251966 555744
rect 226886 555063 226891 555249
rect 227077 555063 227082 555249
rect 226886 555058 227082 555063
rect 149540 554689 149640 554694
rect 149540 554599 149545 554689
rect 149635 554599 149640 554689
rect 149540 554594 149640 554599
rect 136929 553124 142918 553302
rect 142360 553122 142906 553124
rect 135565 552836 142920 553014
rect 142362 552834 142908 552836
rect 134187 552520 142928 552698
rect 142370 552518 142916 552520
rect 180682 552466 227148 552576
rect 132727 552246 142930 552424
rect 180682 552270 226886 552466
rect 227082 552270 227148 552466
rect 142372 552244 142918 552246
rect 131397 551944 142914 552122
rect 180682 552120 227148 552270
rect 142356 551942 142902 551944
rect 130351 551662 142910 551840
rect 142352 551660 142898 551662
rect 129433 551384 142928 551562
rect 142370 551382 142916 551384
rect 128683 551086 142930 551264
rect 142372 551084 142918 551086
rect 14568 550261 74810 550266
rect 14568 550011 14573 550261
rect 14823 550170 74810 550261
rect 14823 550110 74718 550170
rect 74778 550110 74810 550170
rect 14823 550011 74810 550110
rect 14568 550006 74810 550011
rect 7861 549435 149688 549440
rect 7861 549131 7866 549435
rect 8170 549362 149688 549435
rect 8170 549262 149540 549362
rect 149640 549262 149688 549362
rect 8170 549131 149688 549262
rect 7861 549126 149688 549131
rect 7074 548715 150086 548720
rect 7074 548373 7079 548715
rect 7421 548618 150086 548715
rect 7421 548518 149940 548618
rect 150040 548518 150086 548618
rect 7421 548373 150086 548518
rect 7074 548368 150086 548373
rect 9958 547559 102608 547564
rect 9958 547309 9963 547559
rect 10213 547501 102608 547559
rect 10213 547470 102444 547501
rect 10213 547410 82538 547470
rect 82598 547410 102444 547470
rect 10213 547371 102444 547410
rect 102574 547371 102608 547501
rect 10213 547309 102608 547371
rect 9958 547304 102608 547309
rect 22538 544249 92000 544254
rect 22538 543995 22543 544249
rect 22797 544184 92000 544249
rect 22797 544072 91840 544184
rect 91952 544072 92000 544184
rect 22797 543995 92000 544072
rect 22538 543990 92000 543995
rect 90326 541804 90451 541809
rect 29313 541799 90331 541804
rect 29313 541694 29318 541799
rect 29423 541694 90331 541799
rect 29313 541689 90331 541694
rect 90446 541799 93815 541804
rect 90446 541694 93705 541799
rect 93810 541694 93815 541799
rect 90446 541689 93815 541694
rect 90326 541684 90451 541689
rect 180682 539506 181138 552120
rect 182880 551127 324243 551132
rect 182880 551026 323930 551127
rect 182880 550926 182912 551026
rect 183012 550926 323930 551026
rect 182880 550819 323930 550926
rect 324238 550819 324243 551127
rect 182880 550814 324243 550819
rect 225694 548775 326874 548780
rect 225694 548612 326375 548775
rect 225694 548492 225796 548612
rect 225916 548492 326375 548612
rect 225694 548281 326375 548492
rect 326869 548281 326874 548775
rect 225694 548276 326874 548281
rect 26506 539501 181138 539506
rect 26506 539055 26511 539501
rect 26957 539055 181138 539501
rect 26506 539050 181138 539055
rect 20195 537048 20473 537054
rect 20473 536957 396092 537048
rect 20473 536843 395928 536957
rect 396042 536843 396092 536957
rect 20473 536770 396092 536843
rect 20195 536764 20473 536770
rect 21652 536092 22172 536098
rect 22172 535901 322800 536092
rect 22172 535759 322604 535901
rect 322746 535759 322800 535901
rect 22172 535572 322800 535759
rect 21652 535566 22172 535572
rect 22676 534894 23016 534900
rect 23016 534771 249362 534894
rect 23016 534653 249190 534771
rect 249308 534653 249362 534771
rect 23016 534554 249362 534653
rect 22676 534548 23016 534554
rect 29307 534306 29421 534311
rect 19726 534202 29312 534306
rect 29416 534202 29421 534306
rect -800 511530 484 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect 19726 508096 19830 534202
rect 29307 534197 29421 534202
rect 23489 533848 23855 533854
rect 23855 533730 176034 533848
rect 23855 533590 175860 533730
rect 176000 533590 176034 533730
rect 23855 533482 176034 533590
rect 23489 533476 23855 533482
rect 26785 533179 26913 533184
rect 74314 533180 74435 533185
rect 74314 533179 74319 533180
rect 26784 533178 74319 533179
rect 26784 533050 26785 533178
rect 26913 533069 74319 533178
rect 74430 533179 74435 533180
rect 74430 533069 74455 533179
rect 26913 533050 74455 533069
rect 26784 533049 74455 533050
rect 26785 533044 26913 533049
rect 27019 532939 27151 532944
rect 27018 532938 98755 532939
rect 27018 532806 27019 532938
rect 27151 532934 98755 532938
rect 27151 532810 98626 532934
rect 98750 532810 98755 532934
rect 27151 532806 98755 532810
rect 27018 532805 98755 532806
rect 27019 532800 27151 532805
rect 27247 532689 27379 532694
rect 27246 532688 99187 532689
rect 27246 532556 27247 532688
rect 27379 532684 99187 532688
rect 27379 532560 99058 532684
rect 99182 532560 99187 532684
rect 27379 532556 99187 532560
rect 27246 532555 99187 532556
rect 27247 532550 27379 532555
rect 27483 532442 27609 532447
rect 27482 532441 99598 532442
rect 27482 532315 27483 532441
rect 27609 532437 99598 532441
rect 27609 532319 99475 532437
rect 99593 532319 99598 532437
rect 27609 532315 99598 532319
rect 27482 532314 99598 532315
rect 27483 532309 27609 532314
rect 27715 532220 27833 532225
rect 27714 532219 100090 532220
rect 27714 532101 27715 532219
rect 27833 532215 100090 532219
rect 27833 532105 99975 532215
rect 100085 532105 100090 532215
rect 27833 532101 100090 532105
rect 27714 532100 100090 532101
rect 27715 532095 27833 532100
rect 27945 531965 28073 531970
rect 27944 531964 100593 531965
rect 27944 531836 27945 531964
rect 28073 531960 100593 531964
rect 28073 531840 100468 531960
rect 100588 531840 100593 531960
rect 28073 531836 100593 531840
rect 27944 531835 100593 531836
rect 27945 531830 28073 531835
rect 28177 531690 28339 531695
rect 28176 531689 101060 531690
rect 28176 531527 28177 531689
rect 28339 531685 101060 531689
rect 28339 531531 100901 531685
rect 101055 531531 101060 531685
rect 28339 531527 101060 531531
rect 28176 531526 101060 531527
rect 28177 531521 28339 531526
rect 542574 531466 543419 531538
rect 542574 531406 542602 531466
rect 542662 531406 543419 531466
rect 28483 531355 28639 531360
rect 28482 531354 101521 531355
rect 28482 531198 28483 531354
rect 28639 531350 101521 531354
rect 28639 531202 101368 531350
rect 101516 531202 101521 531350
rect 542574 531336 543419 531406
rect 543621 531336 543627 531538
rect 28639 531198 101521 531202
rect 28482 531197 101521 531198
rect 28483 531192 28639 531197
rect 469322 531060 543425 531122
rect 28811 531040 28965 531045
rect 28810 531039 101940 531040
rect 28810 530885 28811 531039
rect 28965 531035 101940 531039
rect 28965 530889 101789 531035
rect 101935 530889 101940 531035
rect 469322 530970 469350 531060
rect 469440 530970 543425 531060
rect 469322 530936 543425 530970
rect 543611 530936 543617 531122
rect 28965 530885 101940 530889
rect 28810 530884 101940 530885
rect 28811 530879 28965 530884
rect 24253 530678 24387 530684
rect 24387 530646 27942 530678
rect 24387 530586 27862 530646
rect 27922 530586 27942 530646
rect 24387 530544 27942 530586
rect 24253 530538 24387 530544
rect -800 507984 19830 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 24593 500484 24711 500490
rect 24711 500454 27734 500484
rect 24711 500394 27658 500454
rect 27718 500394 27734 500454
rect 24711 500366 27734 500394
rect 24593 500360 24711 500366
rect 24913 470292 25031 470298
rect 25031 470262 27734 470292
rect 25031 470202 27658 470262
rect 27718 470202 27734 470262
rect 25031 470174 27734 470202
rect 24913 470168 25031 470174
rect -800 468415 17160 468420
rect -800 468313 17053 468415
rect 17155 468313 17160 468415
rect -800 468308 17160 468313
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 25215 440100 25333 440106
rect 25333 440070 27734 440100
rect 25333 440010 27658 440070
rect 27718 440010 27734 440070
rect 25333 439982 27734 440010
rect 25215 439976 25333 439982
rect -800 425193 22728 425198
rect -800 425091 22621 425193
rect 22723 425091 22728 425193
rect -800 425086 22728 425091
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 25493 409976 25611 409982
rect 25611 409946 27734 409976
rect 25611 409886 27658 409946
rect 27718 409886 27734 409946
rect 25611 409858 27734 409886
rect 25493 409852 25611 409858
rect -800 381971 12344 381976
rect -800 381869 12237 381971
rect 12339 381869 12344 381971
rect -800 381864 12344 381869
rect -800 380682 480 380794
rect 25783 379784 25901 379790
rect 25901 379754 27734 379784
rect 25901 379694 27658 379754
rect 27718 379694 27734 379754
rect 25901 379666 27734 379694
rect 25783 379660 25901 379666
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 26065 349592 26183 349598
rect 26183 349562 27734 349592
rect 26183 349502 27658 349562
rect 27718 349502 27734 349562
rect 26183 349474 27734 349502
rect 26065 349468 26183 349474
rect -800 338749 4710 338754
rect -800 338647 4603 338749
rect 4705 338647 4710 338749
rect -800 338642 4710 338647
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 26317 319468 26435 319474
rect 26435 319438 27734 319468
rect 26435 319378 27658 319438
rect 27718 319378 27734 319438
rect 26435 319350 27734 319378
rect 26317 319344 26435 319350
rect -800 295527 26806 295532
rect -800 295425 26699 295527
rect 26801 295425 26806 295527
rect -800 295420 26806 295425
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect 26554 289694 26674 289700
rect -800 289510 480 289622
rect 26554 289246 26674 289574
rect 26554 289186 26586 289246
rect 26646 289186 26674 289246
rect 26554 289152 26674 289186
rect 544900 269342 547088 582000
rect 550536 313764 552174 587608
rect 552788 530658 553106 530704
rect 552788 530568 552899 530658
rect 552989 530568 553106 530658
rect 552788 530380 553106 530568
rect 552788 530280 552790 530380
rect 552790 530058 553106 530064
rect 556590 358986 558426 611640
rect 563126 405408 563858 617290
rect 568791 449830 569437 621228
rect 573656 494252 574212 623396
rect 577070 583674 577818 627634
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 577070 583562 584800 583674
rect 577070 583558 577818 583562
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 573656 494140 584800 494252
rect 573656 494138 574212 494140
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 568791 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 563126 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 556590 358878 584800 358986
rect 556632 358874 584800 358878
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 550536 313652 584800 313764
rect 583520 275140 584800 275252
rect 555634 274218 555886 274260
rect 555634 274158 555728 274218
rect 555788 274158 555886 274218
rect 555634 273956 555886 274158
rect 583520 273958 584800 274070
rect 555634 273698 555886 273704
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 544900 269230 584800 269342
rect 26784 259296 26914 259302
rect 26784 259054 26914 259166
rect 26784 258994 26818 259054
rect 26878 258994 26914 259054
rect 26784 258976 26914 258994
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248959 14710 248964
rect -800 248857 14603 248959
rect 14705 248857 14710 248959
rect -800 248852 14710 248857
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 27018 229058 27152 229064
rect 27018 228862 27152 228924
rect 27018 228802 27056 228862
rect 27116 228802 27152 228862
rect 27018 228780 27152 228802
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 27246 198980 27380 198986
rect 27246 198738 27380 198846
rect 27246 198678 27284 198738
rect 27344 198678 27380 198738
rect 27246 198662 27380 198678
rect 548619 195130 549289 195135
rect 582340 195130 584800 196230
rect 548618 195129 584800 195130
rect 548618 194459 548619 195129
rect 549289 194459 584800 195129
rect 548618 194458 584800 194459
rect 548619 194453 549289 194458
rect 548673 184250 549343 184255
rect 577294 184250 577966 194458
rect 582340 191430 584800 194458
rect 582340 184250 584800 186230
rect 548672 184249 584800 184250
rect 548672 183579 548673 184249
rect 549343 183579 584800 184249
rect 548672 183578 584800 183579
rect 548673 183573 549343 183578
rect 582340 181430 584800 183578
rect -800 172888 1660 177688
rect 27482 168746 27610 168752
rect 27482 168546 27610 168618
rect 27482 168486 27518 168546
rect 27578 168486 27610 168546
rect 27482 168466 27610 168486
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 27714 138568 27834 138574
rect 27714 138354 27834 138448
rect 27714 138294 27752 138354
rect 27812 138294 27834 138354
rect 27714 138278 27834 138294
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121337 10102 121342
rect -800 121235 9995 121337
rect 10097 121235 10102 121337
rect -800 121230 10102 121235
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 27944 108478 28074 108484
rect 27944 108230 28074 108348
rect 27944 108170 27976 108230
rect 28036 108170 28074 108230
rect 27944 108146 28074 108170
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 580272 92861 584800 92866
rect 580272 92759 580277 92861
rect 580379 92759 584800 92861
rect 580272 92754 584800 92759
rect 583520 91572 584800 91684
rect -800 81661 7272 81666
rect -800 81559 7165 81661
rect 7267 81559 7272 81661
rect -800 81554 7272 81559
rect -800 80372 480 80484
rect -800 79190 480 79302
rect 28176 78516 28340 78522
rect -800 78008 480 78120
rect 28176 78038 28340 78352
rect 28176 77978 28230 78038
rect 28290 77978 28340 78038
rect 28176 77950 28340 77978
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 567598 48203 584800 48208
rect 567598 48101 567603 48203
rect 567705 48101 584800 48203
rect 567598 48096 584800 48101
rect 28482 48072 28640 48078
rect 28482 47846 28640 47914
rect 28482 47786 28522 47846
rect 28582 47786 28640 47846
rect 28482 47752 28640 47786
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect 23608 34898 23720 34904
rect -800 34786 23608 34898
rect 23608 34780 23720 34786
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 547614 21750 547726 21756
rect 547726 21638 584800 21750
rect 547614 21632 547726 21638
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 28810 18020 28966 18026
rect 28810 17722 28966 17864
rect 28810 17662 28864 17722
rect 28924 17662 28966 17722
rect 28810 17642 28966 17662
rect 558896 17722 559126 17742
rect 558896 17662 558978 17722
rect 559038 17662 559126 17722
rect 558896 17574 559126 17662
rect 558896 17338 559126 17344
rect 549942 17022 550054 17028
rect -800 16910 480 17022
rect 550054 16910 584800 17022
rect 549942 16904 550054 16910
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect 535055 14918 535725 14923
rect 535054 14917 578558 14918
rect -800 14546 480 14658
rect 535054 14247 535055 14917
rect 535725 14662 578558 14917
rect 535725 14540 578199 14662
rect 578321 14540 578558 14662
rect 582044 14653 584800 14658
rect 582044 14551 582049 14653
rect 582151 14551 584800 14653
rect 582044 14546 584800 14551
rect 535725 14247 578558 14540
rect 535054 14246 578558 14247
rect 535055 14241 535725 14246
rect 22804 13476 22916 13482
rect -800 13364 22804 13476
rect 22804 13358 22916 13364
rect 552908 13476 553020 13482
rect 553020 13364 584800 13476
rect 552908 13358 553020 13364
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect 582056 9930 583806 9932
rect -800 9818 480 9930
rect 582056 9927 584800 9930
rect 582056 9825 582061 9927
rect 582163 9825 584800 9927
rect 582056 9820 584800 9825
rect 583520 9818 584800 9820
rect 21858 8748 21970 8754
rect -800 8636 21858 8748
rect 21858 8630 21970 8636
rect 555718 8748 555830 8754
rect 555830 8636 584800 8748
rect 555718 8630 555830 8636
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 582168 5197 584800 5202
rect 582168 5095 582173 5197
rect 582275 5095 584800 5197
rect 582168 5090 584800 5095
rect 20274 4020 20386 4026
rect -800 3908 20274 4020
rect 20274 3902 20386 3908
rect 558952 4020 559064 4026
rect 559064 3908 584800 4020
rect 558952 3902 559064 3908
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 412641 698770 413247 699376
rect 30406 689916 34854 690814
rect 417384 699249 417736 699254
rect 417384 698912 417389 699249
rect 417389 698912 417731 699249
rect 417731 698912 417736 699249
rect 470540 699255 470904 699260
rect 470540 698906 470545 699255
rect 470545 698906 470899 699255
rect 470899 698906 470904 699255
rect 520568 696744 523028 699204
rect 512816 692626 515276 695086
rect 560023 689712 560397 689717
rect 560023 689353 560028 689712
rect 560028 689353 560392 689712
rect 560392 689353 560397 689712
rect 15002 643900 19666 648564
rect 575938 639830 580658 644550
rect 137841 620281 137991 620431
rect 140292 620282 140440 620430
rect 24254 594432 24386 594564
rect 24594 594146 24710 594262
rect 24914 593850 25030 593966
rect 25216 593582 25332 593698
rect 25494 593312 25610 593428
rect 25784 593000 25900 593116
rect 26066 592710 26182 592826
rect 26318 592420 26434 592536
rect 26555 592149 26673 592267
rect 20195 536770 20473 537048
rect 21652 535572 22172 536092
rect 22676 534554 23016 534894
rect 23489 533482 23855 533848
rect 26785 533050 26913 533178
rect 27019 532806 27151 532938
rect 27247 532556 27379 532688
rect 27483 532315 27609 532441
rect 27715 532101 27833 532219
rect 27945 531836 28073 531964
rect 28177 531527 28339 531689
rect 28483 531198 28639 531354
rect 543419 531336 543621 531538
rect 28811 530885 28965 531039
rect 543425 530936 543611 531122
rect 24253 530544 24387 530678
rect 24593 500366 24711 500484
rect 24913 470174 25031 470292
rect 25215 439982 25333 440100
rect 25493 409858 25611 409976
rect 25783 379666 25901 379784
rect 26065 349474 26183 349592
rect 26317 319350 26435 319468
rect 26554 289574 26674 289694
rect 552790 530064 553106 530380
rect 555634 273704 555886 273956
rect 26784 259166 26914 259296
rect 27018 228924 27152 229058
rect 27246 198846 27380 198980
rect 548619 194459 549289 195129
rect 548673 183579 549343 184249
rect 27482 168618 27610 168746
rect 27714 138448 27834 138568
rect 27944 108348 28074 108478
rect 28176 78352 28340 78516
rect 28482 47914 28640 48072
rect 23608 34786 23720 34898
rect 547614 21638 547726 21750
rect 28810 17864 28966 18020
rect 558896 17344 559126 17574
rect 549942 16910 550054 17022
rect 535055 14247 535725 14917
rect 22804 13364 22916 13476
rect 552908 13364 553020 13476
rect 21858 8636 21970 8748
rect 555718 8636 555830 8748
rect 20274 3908 20386 4020
rect 558952 3908 559064 4020
<< metal4 >>
rect 412640 699376 413248 699377
rect 412640 698770 412641 699376
rect 413247 699260 561426 699376
rect 413247 699254 470540 699260
rect 413247 698912 417384 699254
rect 417736 698912 470540 699254
rect 413247 698906 470540 698912
rect 470904 699204 561426 699260
rect 470904 698906 520568 699204
rect 413247 698770 520568 698906
rect 412640 698769 413248 698770
rect 505280 696744 520568 698770
rect 523028 696744 561436 699204
rect 520567 696743 523029 696744
rect 512815 695086 515277 695087
rect 512815 692626 512816 695086
rect 515276 692626 515277 695086
rect 512815 692625 515277 692626
rect 30276 690814 34940 691006
rect 30276 689916 30406 690814
rect 34854 689916 34940 690814
rect 15001 648564 19667 648565
rect 30276 648564 34940 689916
rect 512816 677318 515276 692625
rect 558976 689717 561436 696744
rect 558976 689353 560023 689717
rect 560397 689353 561436 689717
rect 558976 689304 561436 689353
rect 335440 665430 515346 677318
rect 15001 643900 15002 648564
rect 19666 646916 79422 648564
rect 19666 643900 79482 646916
rect 15001 643899 19667 643900
rect 77850 641872 79482 643900
rect 77850 641072 101504 641872
rect 77850 641066 79482 641072
rect 85622 641066 87254 641072
rect 335440 633052 347328 665430
rect 575937 644550 580659 644551
rect 537992 644546 575938 644550
rect 319632 632252 347328 633052
rect 335440 632248 347328 632252
rect 535732 639830 575938 644546
rect 580658 639830 580659 644550
rect 77850 618834 79482 620798
rect 85622 618834 87254 620798
rect 137840 620431 137992 620432
rect 137840 620281 137841 620431
rect 137991 620430 140441 620431
rect 137991 620282 140292 620430
rect 140440 620282 140441 620430
rect 137991 620281 140441 620282
rect 137840 620280 137992 620281
rect 24253 594564 24387 594565
rect 24253 594432 24254 594564
rect 24386 594432 24387 594564
rect 20194 537048 20474 537049
rect 20194 536770 20195 537048
rect 20473 536770 20474 537048
rect 20194 536769 20474 536770
rect 20195 4020 20473 536769
rect 21651 536092 22173 536093
rect 21651 535572 21652 536092
rect 22172 535572 22173 536092
rect 21651 535571 22173 535572
rect 21652 8748 22172 535571
rect 22675 534894 23017 534895
rect 22675 534554 22676 534894
rect 23016 534554 23017 534894
rect 22675 534553 23017 534554
rect 22676 13476 23016 534553
rect 23488 533848 23856 533849
rect 23488 533482 23489 533848
rect 23855 533482 23856 533848
rect 23488 533481 23856 533482
rect 23489 34898 23855 533481
rect 24253 530679 24387 594432
rect 24593 594262 24711 594263
rect 24593 594146 24594 594262
rect 24710 594146 24711 594262
rect 24252 530678 24388 530679
rect 24252 530544 24253 530678
rect 24387 530544 24388 530678
rect 24252 530543 24388 530544
rect 24593 500485 24711 594146
rect 24913 593966 25031 593967
rect 24913 593850 24914 593966
rect 25030 593850 25031 593966
rect 24592 500484 24712 500485
rect 24592 500366 24593 500484
rect 24711 500366 24712 500484
rect 24592 500365 24712 500366
rect 24913 470293 25031 593850
rect 25215 593698 25333 593699
rect 25215 593582 25216 593698
rect 25332 593582 25333 593698
rect 24912 470292 25032 470293
rect 24912 470174 24913 470292
rect 25031 470174 25032 470292
rect 24912 470173 25032 470174
rect 25215 440101 25333 593582
rect 25493 593428 25611 593429
rect 25493 593312 25494 593428
rect 25610 593312 25611 593428
rect 25214 440100 25334 440101
rect 25214 439982 25215 440100
rect 25333 439982 25334 440100
rect 25214 439981 25334 439982
rect 25493 409977 25611 593312
rect 25783 593116 25901 593117
rect 25783 593000 25784 593116
rect 25900 593000 25901 593116
rect 25492 409976 25612 409977
rect 25492 409858 25493 409976
rect 25611 409858 25612 409976
rect 25492 409857 25612 409858
rect 25783 379785 25901 593000
rect 26065 592826 26183 592827
rect 26065 592710 26066 592826
rect 26182 592710 26183 592826
rect 25782 379784 25902 379785
rect 25782 379666 25783 379784
rect 25901 379666 25902 379784
rect 25782 379665 25902 379666
rect 26065 349593 26183 592710
rect 26317 592536 26435 592537
rect 26317 592420 26318 592536
rect 26434 592420 26435 592536
rect 26064 349592 26184 349593
rect 26064 349474 26065 349592
rect 26183 349474 26184 349592
rect 26064 349473 26184 349474
rect 26317 319469 26435 592420
rect 26554 592267 26674 592268
rect 26554 592149 26555 592267
rect 26673 592149 26674 592267
rect 26316 319468 26436 319469
rect 26316 319350 26317 319468
rect 26435 319350 26436 319468
rect 26316 319349 26436 319350
rect 26554 289695 26674 592149
rect 75402 566818 77034 607942
rect 77850 600360 79482 605350
rect 85622 600360 87254 605302
rect 77848 599560 87254 600360
rect 77850 567218 79482 599560
rect 85622 568074 87254 599560
rect 88070 568472 89702 607942
rect 75418 534000 77050 556592
rect 77866 549010 79498 554000
rect 85638 549010 87270 553952
rect 77864 548210 87270 549010
rect 26784 533178 26914 533179
rect 26784 533050 26785 533178
rect 26913 533050 26914 533178
rect 26553 289694 26675 289695
rect 26553 289574 26554 289694
rect 26674 289574 26675 289694
rect 26553 289573 26675 289574
rect 26784 259297 26914 533050
rect 27018 532938 27152 532939
rect 27018 532806 27019 532938
rect 27151 532806 27152 532938
rect 26783 259296 26915 259297
rect 26783 259166 26784 259296
rect 26914 259166 26915 259296
rect 26783 259165 26915 259166
rect 27018 229059 27152 532806
rect 27246 532688 27380 532689
rect 27246 532556 27247 532688
rect 27379 532556 27380 532688
rect 27017 229058 27153 229059
rect 27017 228924 27018 229058
rect 27152 228924 27153 229058
rect 27017 228923 27153 228924
rect 27246 198981 27380 532556
rect 27482 532441 27610 532442
rect 27482 532315 27483 532441
rect 27609 532315 27610 532441
rect 75418 532368 78776 534000
rect 27245 198980 27381 198981
rect 27245 198846 27246 198980
rect 27380 198846 27381 198980
rect 27245 198845 27381 198846
rect 27482 168747 27610 532315
rect 27714 532219 27834 532220
rect 27714 532101 27715 532219
rect 27833 532101 27834 532219
rect 27481 168746 27611 168747
rect 27481 168618 27482 168746
rect 27610 168618 27611 168746
rect 27481 168617 27611 168618
rect 27714 138569 27834 532101
rect 27944 531964 28074 531965
rect 27944 531836 27945 531964
rect 28073 531836 28074 531964
rect 27713 138568 27835 138569
rect 27713 138448 27714 138568
rect 27834 138448 27835 138568
rect 27713 138447 27835 138448
rect 27944 108479 28074 531836
rect 28176 531689 28340 531690
rect 28176 531527 28177 531689
rect 28339 531527 28340 531689
rect 27943 108478 28075 108479
rect 27943 108348 27944 108478
rect 28074 108348 28075 108478
rect 27943 108347 28075 108348
rect 28176 78517 28340 531527
rect 28482 531354 28640 531355
rect 28482 531198 28483 531354
rect 28639 531198 28640 531354
rect 28175 78516 28341 78517
rect 28175 78352 28176 78516
rect 28340 78352 28341 78516
rect 28175 78351 28341 78352
rect 28482 48073 28640 531198
rect 28810 531039 28966 531040
rect 28810 530885 28811 531039
rect 28965 530885 28966 531039
rect 28481 48072 28641 48073
rect 28481 47914 28482 48072
rect 28640 47914 28641 48072
rect 28481 47913 28641 47914
rect 23489 34786 23608 34898
rect 23720 34786 23855 34898
rect 23489 34720 23855 34786
rect 28810 18021 28966 530885
rect 78094 500366 78766 532368
rect 80746 531852 81546 548210
rect 88086 532276 89718 554700
rect 535732 532446 541064 639830
rect 575937 639829 580659 639830
rect 80814 496902 81486 531852
rect 88974 504554 89646 532276
rect 537882 510238 539514 532446
rect 543418 531538 543622 531539
rect 543418 531336 543419 531538
rect 543621 531336 550107 531538
rect 543418 531335 543622 531336
rect 543424 531122 543612 531123
rect 543424 530936 543425 531122
rect 543611 530936 547764 531122
rect 543424 530935 543612 530936
rect 28809 18020 28967 18021
rect 28809 17864 28810 18020
rect 28966 17864 28967 18020
rect 28809 17863 28967 17864
rect 535054 14917 535726 39862
rect 547578 21750 547764 530936
rect 548618 195129 549290 195130
rect 548618 194459 548619 195129
rect 549289 194459 549290 195129
rect 548618 194458 549290 194459
rect 548672 184249 549344 184250
rect 548672 183579 548673 184249
rect 549343 183579 549344 184249
rect 548672 183578 549344 183579
rect 547578 21638 547614 21750
rect 547726 21638 547764 21750
rect 547578 21599 547764 21638
rect 549905 17022 550107 531336
rect 552789 530380 553107 530381
rect 549905 16910 549942 17022
rect 550054 16910 550107 17022
rect 549905 16879 550107 16910
rect 552784 530064 552790 530380
rect 553106 530206 553110 530380
rect 553106 530064 553112 530206
rect 535054 14247 535055 14917
rect 535725 14247 535726 14917
rect 535054 14246 535726 14247
rect 22676 13364 22804 13476
rect 22916 13364 23016 13476
rect 22676 13346 23016 13364
rect 552784 13476 553112 530064
rect 555633 273956 555887 273957
rect 555633 273704 555634 273956
rect 555886 273704 555887 273956
rect 555633 273703 555887 273704
rect 552784 13364 552908 13476
rect 553020 13364 553112 13476
rect 552784 13322 553112 13364
rect 21652 8636 21858 8748
rect 21970 8636 22172 8748
rect 21652 8596 22172 8636
rect 555634 8748 555886 273703
rect 558895 17574 559127 17575
rect 558895 17344 558896 17574
rect 559126 17344 559127 17574
rect 558895 17343 559127 17344
rect 555634 8636 555718 8748
rect 555830 8636 555886 8748
rect 555634 8596 555886 8636
rect 20195 3908 20274 4020
rect 20386 3908 20473 4020
rect 20195 3871 20473 3908
rect 558896 4020 559126 17343
rect 558896 3908 558952 4020
rect 559064 3908 559126 4020
rect 558896 3869 559126 3908
<< via4 >>
rect 548642 194482 549266 195106
rect 548696 183602 549320 184226
<< metal5 >>
rect 93520 621340 93548 621350
rect 539778 195106 549290 195130
rect 539778 194482 548642 195106
rect 549266 194482 549290 195106
rect 539778 194458 549290 194482
rect 540754 184226 549344 184250
rect 540754 183602 548696 184226
rect 549320 183602 549344 184226
rect 540754 183578 549344 183602
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_0
timestamp 1624477805
transform 0 1 579723 -1 0 5146
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_1
timestamp 1624477805
transform 0 1 579611 -1 0 9876
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_2
timestamp 1624477805
transform 0 1 579599 -1 0 14602
box -60 -357 60 357
use sar_adc_controller_8bit  sar_adc_controller_8bit_0
timestamp 1624477805
transform -1 0 90618 0 -1 570806
box 0 0 16100 20128
use sar_adc_controller_8bit  sar_adc_controller_8bit_1
timestamp 1624477805
transform -1 0 90602 0 -1 622156
box 0 0 16100 20128
use analog_top_level  analog_top_level_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/analog_top_level
timestamp 1624477805
transform -1 0 479200 0 1 739592
box 157324 -188462 385680 -59028
use esd_cell  esd_cell_1 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/esd_cell
timestamp 1624477805
transform 1 0 5996 0 1 682782
box -2400 -3178 2400 3178
use esd_cell  esd_cell_0
timestamp 1624477805
transform 1 0 22248 0 1 697476
box -2400 -3178 2400 3178
use esd_cell  esd_cell_2
timestamp 1624477805
transform 1 0 75404 0 1 697476
box -2400 -3178 2400 3178
use esd_cell  esd_cell_3
timestamp 1624477805
transform 1 0 127332 0 1 698616
box -2400 -3178 2400 3178
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_4
timestamp 1624477805
transform -1 0 174470 0 -1 701565
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_3
timestamp 1624477805
transform -1 0 171964 0 -1 701565
box -60 -357 60 357
use esd_cell  esd_cell_5
timestamp 1624477805
transform 1 0 215186 0 1 695212
box -2400 -3178 2400 3178
use esd_cell  esd_cell_4
timestamp 1624477805
transform 1 0 200032 0 1 689638
box -2400 -3178 2400 3178
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_5
timestamp 1624477805
transform -1 0 223752 0 -1 701565
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_6
timestamp 1624477805
transform -1 0 226152 0 -1 701565
box -60 -357 60 357
use esd_cell  esd_cell_7
timestamp 1624477805
transform 1 0 408838 0 1 696756
box -2400 -3178 2400 3178
use esd_cell  esd_cell_6
timestamp 1624477805
transform 1 0 318206 0 1 694824
box -2400 -3178 2400 3178
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_8
timestamp 1624477805
transform -1 0 327900 0 -1 701565
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_7
timestamp 1624477805
transform -1 0 325390 0 -1 701565
box -60 -357 60 357
use esd_cell  esd_cell_8
timestamp 1624477805
transform 1 0 463684 0 1 693044
box -2400 -3178 2400 3178
use esd_cell  esd_cell_10
timestamp 1624477805
transform 1 0 577108 0 1 680432
box -2400 -3178 2400 3178
use esd_cell  esd_cell_9
timestamp 1624477805
transform 1 0 566444 0 1 692528
box -2400 -3178 2400 3178
use deconv_kernel_estimator_top_level  deconv_kernel_estimator_top_level_0
timestamp 1624477805
transform 1 0 29134 0 1 17658
box 0 0 513728 512992
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1400 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1400 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1400 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1400 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1400 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1400 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1400 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1400 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1400 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1400 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1400 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1400 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1400 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1400 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1400 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1400 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1400 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1400 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1400 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1400 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1400 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1400 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1400 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1400 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1400 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1400 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1400 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1400 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1400 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1400 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1400 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1400 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1400 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1400 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 2400 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 2400 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 2400 180 0 0 io_analog[3]
port 41 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 2400 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 2400 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 2400 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 2400 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 2400 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 2400 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 2400 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1400 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1400 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1400 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1400 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1400 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1400 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1400 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1400 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1400 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1400 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1400 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1400 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1400 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1400 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1400 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1400 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1400 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1400 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1400 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1400 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1400 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1400 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1400 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1400 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1400 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1400 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1400 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1400 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1400 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1400 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1400 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1400 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1400 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1400 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1400 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1400 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1400 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1400 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1400 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1400 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1400 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1400 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1400 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1400 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1400 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1400 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1400 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1400 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1400 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1400 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1400 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1400 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1400 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1400 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1400 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1400 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1400 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1400 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1400 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1400 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1400 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1400 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1400 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1400 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1400 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1400 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1400 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1400 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1400 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1400 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1400 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1400 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1400 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1400 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1400 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1400 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1400 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1400 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1400 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1400 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1400 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1400 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1400 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1400 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1400 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1400 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1400 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1400 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1400 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1400 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1400 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1400 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1400 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1400 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1400 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1400 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1400 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1400 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1400 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1400 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1400 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1400 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1400 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1400 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1400 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1400 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1400 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1400 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1400 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1400 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1400 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1400 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1400 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1400 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1400 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1400 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1400 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1400 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1400 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1400 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1400 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1400 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1400 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1400 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1400 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1400 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1400 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1400 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1400 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1400 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1400 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1400 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1400 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1400 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1400 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1400 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1400 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1400 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1400 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1400 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1400 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1400 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1400 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1400 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1400 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1400 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1400 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1400 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1400 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1400 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1400 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1400 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1400 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1400 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1400 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1400 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1400 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1400 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1400 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1400 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1400 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1400 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1400 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1400 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1400 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1400 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1400 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1400 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1400 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1400 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1400 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1400 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1400 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1400 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1400 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1400 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1400 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1400 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1400 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1400 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1400 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1400 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1400 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1400 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1400 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1400 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1400 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1400 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1400 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1400 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1400 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1400 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1400 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1400 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1400 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1400 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1400 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1400 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1400 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1400 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1400 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1400 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1400 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1400 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1400 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1400 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1400 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1400 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1400 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1400 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1400 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1400 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1400 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1400 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1400 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1400 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1400 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1400 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1400 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1400 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1400 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1400 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1400 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1400 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1400 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1400 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1400 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1400 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1400 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1400 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1400 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1400 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1400 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1400 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1400 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1400 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1400 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1400 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1400 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1400 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1400 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1400 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1400 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1400 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1400 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1400 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1400 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1400 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1400 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1400 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1400 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1400 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1400 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1400 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1400 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1400 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1400 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1400 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1400 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1400 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1400 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1400 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1400 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1400 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1400 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1400 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1400 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1400 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1400 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1400 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1400 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1400 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1400 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1400 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1400 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1400 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1400 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1400 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1400 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1400 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1400 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1400 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1400 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1400 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1400 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1400 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1400 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1400 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1400 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1400 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1400 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1400 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1400 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1400 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1400 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1400 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1400 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1400 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1400 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1400 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1400 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1400 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1400 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1400 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1400 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1400 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1400 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1400 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1400 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1400 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1400 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1400 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1400 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1400 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1400 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1400 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1400 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1400 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1400 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1400 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1400 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1400 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1400 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1400 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1400 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1400 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1400 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1400 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1400 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1400 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1400 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1400 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1400 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1400 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1400 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1400 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1400 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1400 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1400 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1400 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1400 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1400 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1400 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1400 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1400 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1400 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1400 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1400 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1400 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1400 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1400 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1400 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1400 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1400 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1400 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1400 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1400 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1400 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1400 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1400 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1400 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1400 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1400 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1400 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1400 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1400 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1400 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1400 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1400 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1400 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1400 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1400 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1400 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1400 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1400 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1400 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1400 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1400 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1400 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1400 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1400 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1400 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1400 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1400 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1400 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1400 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1400 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1400 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1400 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1400 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1400 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1400 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1400 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1400 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1400 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1400 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1400 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1400 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1400 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1400 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1400 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1400 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1400 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1400 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1400 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1400 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1400 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1400 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1400 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1400 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1400 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1400 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1400 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1400 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1400 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1400 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1400 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1400 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1400 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1400 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1400 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1400 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1400 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1400 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1400 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1400 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1400 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1400 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1400 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1400 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1400 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1400 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1400 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1400 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1400 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1400 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1400 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1400 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1400 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1400 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1400 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1400 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1400 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1400 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1400 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1400 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1400 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1400 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1400 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1400 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1400 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1400 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1400 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1400 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1400 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1400 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1400 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1400 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1400 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1400 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1400 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1400 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1400 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1400 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1400 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1400 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1400 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1400 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1400 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1400 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1400 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1400 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1400 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1400 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1400 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1400 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1400 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1400 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1400 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1400 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1400 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1400 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1400 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1400 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1400 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1400 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1400 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1400 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1400 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1400 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1400 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1400 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1400 0 0 0 vdda2
port 553 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1400 0 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1400 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1400 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1400 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1400 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1400 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1400 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1400 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1400 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1400 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1400 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1400 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1400 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1400 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1400 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1400 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1400 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1400 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1400 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1400 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1400 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1400 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1400 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1400 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1400 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1400 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1400 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1400 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1400 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1400 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1400 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1400 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1400 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1400 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1400 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1400 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1400 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1400 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1400 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1400 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1400 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1400 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1400 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1400 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1400 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1400 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1400 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1400 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1400 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1400 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1400 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1400 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1400 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1400 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1400 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1400 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1400 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1400 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1400 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1400 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1400 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1400 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1400 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1400 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1400 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1400 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1400 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1400 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1400 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1400 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1400 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1400 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1400 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1400 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1400 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1400 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1400 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1400 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1400 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1400 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1400 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1400 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1400 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1400 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1400 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1400 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1400 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1400 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1400 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1400 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1400 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1400 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1400 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1400 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1400 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1400 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1400 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1400 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1400 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1400 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1400 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1400 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1400 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1400 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1400 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1400 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1400 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1400 90 0 0 wbs_we_i
port 663 nsew
flabel metal3 97138 619918 97180 619954 1 FreeSans 480 0 0 0 sig_frequency_7
flabel metal3 97036 617672 97078 617714 1 FreeSans 480 0 0 0 sig_frequency_6
flabel metal3 96998 615414 97028 615456 1 FreeSans 480 0 0 0 sig_frequency_5
flabel metal3 96882 613170 96918 613214 1 FreeSans 480 0 0 0 sig_frequency_4
flabel metal3 96900 610990 96924 611028 1 FreeSans 480 0 0 0 sig_frequency_3
flabel metal3 96764 608770 96790 608796 1 FreeSans 480 0 0 0 sig_frequency_2
flabel metal3 96722 606516 96752 606564 1 FreeSans 480 0 0 0 sig_frequency_1
flabel metal3 96746 604278 96802 604328 1 FreeSans 480 0 0 0 sig_frequency_0
flabel metal3 137200 620356 137222 620376 1 FreeSans 480 0 0 0 sample
flabel metal3 97254 552942 97336 552992 1 FreeSans 480 0 0 0 sig_amplitude_0
flabel metal3 97126 555166 97172 555212 1 FreeSans 480 0 0 0 sig_amplitude_1
flabel metal3 96984 557436 97020 557470 1 FreeSans 480 0 0 0 sig_amplitude_2
flabel metal3 96762 559642 96798 559674 1 FreeSans 480 0 0 0 sig_amplitude_3
flabel metal3 96656 561850 96696 561878 1 FreeSans 480 0 0 0 sig_amplitude_4
flabel metal3 96516 564072 96548 564108 1 FreeSans 480 0 0 0 sig_amplitude_5
flabel metal3 96390 566330 96434 566374 1 FreeSans 480 0 0 0 sig_amplitude_6
flabel metal3 96328 567996 96364 568042 1 FreeSans 480 0 0 0 sig_amplitude_7
flabel metal2 92812 587564 92830 587588 1 FreeSans 480 0 0 0 amplitude_comparator_val
flabel metal2 92824 638576 92846 638598 1 FreeSans 480 0 0 0 frequency_comparator_val
flabel metal3 s -800 511530 480 511642 0 FreeSans 1400 0 0 0 gpio_analog[7]
port 16 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nwell >>
rect 402 846 2798 3698
rect 10 522 2798 846
<< pwell >>
rect 90 214 2798 358
rect 402 -1758 2798 214
<< psubdiff >>
rect 438 222 600 322
rect 2600 222 2762 322
rect 438 160 538 222
rect 438 -1622 538 -1560
rect 2662 160 2762 222
rect 2662 -1622 2762 -1560
rect 438 -1722 600 -1622
rect 2600 -1722 2762 -1622
<< nsubdiff >>
rect 438 3562 600 3662
rect 2600 3562 2762 3662
rect 438 3500 538 3562
rect 438 658 538 720
rect 2662 3500 2762 3562
rect 2662 658 2762 720
rect 438 558 600 658
rect 2600 558 2762 658
<< psubdiffcont >>
rect 600 222 2600 322
rect 438 -1560 538 160
rect 2662 -1560 2762 160
rect 600 -1722 2600 -1622
<< nsubdiffcont >>
rect 600 3562 2600 3662
rect 438 720 538 3500
rect 2662 720 2762 3500
rect 600 558 2600 658
<< locali >>
rect 438 3500 538 3662
rect 438 558 538 720
rect 2662 3500 2762 3662
rect 2662 558 2762 720
rect 438 160 538 322
rect 438 -1722 538 -1560
rect 2662 160 2762 322
rect 2662 -1722 2762 -1560
<< viali >>
rect 538 3562 600 3662
rect 600 3562 2600 3662
rect 2600 3562 2662 3662
rect 438 798 538 3422
rect 2662 798 2762 3422
rect 538 558 600 658
rect 600 558 2600 658
rect 2600 558 2662 658
rect 118 478 166 526
rect 220 420 268 468
rect 538 222 600 322
rect 600 222 2600 322
rect 2600 222 2662 322
rect 438 -1530 538 130
rect 2662 -1530 2762 130
rect 538 -1722 600 -1622
rect 600 -1722 2600 -1622
rect 2600 -1722 2662 -1622
<< metal1 >>
rect 432 3662 2768 3668
rect 432 3562 538 3662
rect 2662 3562 2768 3662
rect 432 3556 2768 3562
rect 432 3422 544 3556
rect 432 854 438 3422
rect 310 798 438 854
rect 538 798 544 3422
rect 1144 3256 1154 3556
rect 2046 3256 2056 3556
rect 2656 3422 2768 3556
rect 700 3052 2602 3082
rect 700 2988 734 3052
rect 2558 2988 2602 3052
rect 700 2958 2602 2988
rect 774 2694 834 2958
rect 904 2694 964 2958
rect 1282 2814 1288 2874
rect 1348 2814 1354 2874
rect 1800 2814 1806 2874
rect 1866 2814 1872 2874
rect 620 2582 626 2642
rect 686 2582 692 2642
rect 774 2634 964 2694
rect 626 2048 686 2582
rect 774 2418 834 2634
rect 904 2506 964 2634
rect 626 1068 686 1988
rect 774 1852 834 2118
rect 904 1852 964 2016
rect 774 1792 964 1852
rect 1030 1804 1090 2100
rect 1160 1918 1220 2016
rect 1154 1858 1160 1918
rect 1220 1858 1226 1918
rect 774 1538 834 1792
rect 904 1648 964 1792
rect 1024 1744 1030 1804
rect 1090 1744 1096 1804
rect 626 1008 876 1068
rect 936 1008 942 1068
rect 1028 956 1088 1260
rect 1288 1252 1348 2814
rect 1538 2702 1544 2762
rect 1604 2702 1610 2762
rect 1410 2582 1416 2642
rect 1476 2582 1482 2642
rect 1416 2506 1476 2582
rect 1544 2418 1604 2702
rect 1666 2582 1672 2642
rect 1732 2582 1738 2642
rect 1672 2504 1732 2582
rect 1806 2390 1866 2814
rect 2194 2682 2254 2958
rect 2322 2682 2382 2958
rect 2468 2702 2474 2762
rect 2534 2702 2540 2762
rect 2194 2622 2382 2682
rect 2194 2508 2254 2622
rect 1412 1858 1418 1918
rect 1478 1858 1484 1918
rect 1670 1858 1676 1918
rect 1736 1858 1742 1918
rect 1418 1650 1478 1858
rect 1542 1744 1548 1804
rect 1608 1744 1614 1804
rect 1548 1558 1608 1744
rect 1676 1654 1736 1858
rect 1800 1546 1860 2132
rect 1934 1918 1994 2016
rect 1928 1858 1934 1918
rect 1994 1858 2000 1918
rect 2064 1804 2124 2124
rect 2322 1860 2382 2622
rect 2058 1744 2064 1804
rect 2124 1744 2130 1804
rect 2190 1800 2382 1860
rect 2190 1650 2250 1800
rect 1160 1068 1220 1158
rect 1154 1008 1160 1068
rect 1220 1008 1226 1068
rect 1022 896 1028 956
rect 1088 896 1094 956
rect 1544 808 1604 1254
rect 1672 1062 1732 1156
rect 1802 848 1862 1268
rect 1936 1068 1996 1160
rect 1930 1008 1936 1068
rect 1996 1008 2002 1068
rect 2064 956 2124 1292
rect 2188 1070 2248 1152
rect 2322 1070 2382 1800
rect 2188 1010 2382 1070
rect 2058 896 2064 956
rect 2124 896 2130 956
rect 310 758 544 798
rect 432 664 544 758
rect 1538 748 1544 808
rect 1604 748 1610 808
rect 1796 788 1802 848
rect 1862 788 1868 848
rect 2188 664 2248 1010
rect 2322 664 2382 1010
rect 2474 956 2534 2702
rect 2468 896 2474 956
rect 2534 896 2540 956
rect 2656 798 2662 3422
rect 2762 798 2768 3422
rect 2656 664 2768 798
rect 432 658 2768 664
rect 432 558 538 658
rect 2662 558 2768 658
rect 432 552 2768 558
rect -108 532 -48 538
rect -48 526 178 532
rect -48 478 118 526
rect 166 478 178 526
rect -48 472 178 478
rect 214 474 274 480
rect -108 466 -48 472
rect 208 414 214 474
rect 274 414 280 474
rect 214 408 274 414
rect 432 322 2768 328
rect 432 310 538 322
rect 314 222 538 310
rect 2662 222 2768 322
rect 314 216 2768 222
rect 314 214 544 216
rect 432 130 544 214
rect 432 -1530 438 130
rect 538 -1530 544 130
rect 1544 168 1604 174
rect 1022 42 1028 102
rect 1088 42 1094 102
rect 1028 -312 1088 42
rect 1276 -2 1282 58
rect 1342 -2 1348 58
rect 1282 -278 1342 -2
rect 1408 -114 1414 -54
rect 1474 -114 1480 -54
rect 1414 -194 1474 -114
rect 1544 -274 1604 108
rect 2656 130 2768 216
rect 1796 -2 1802 58
rect 1862 -2 1868 58
rect 1664 -114 1670 -54
rect 1730 -114 1736 -54
rect 1670 -192 1730 -114
rect 1802 -284 1862 -2
rect 766 -738 826 -564
rect 896 -738 956 -668
rect 766 -798 956 -738
rect 766 -1034 826 -798
rect 896 -1034 956 -798
rect 1022 -864 1082 -582
rect 1156 -750 1216 -666
rect 1930 -750 1990 -666
rect 1150 -810 1156 -750
rect 1216 -810 1222 -750
rect 1924 -810 1930 -750
rect 1990 -810 1996 -750
rect 2058 -864 2118 -564
rect 2186 -744 2246 -668
rect 2314 -744 2374 -572
rect 2186 -804 2374 -744
rect 1016 -924 1022 -864
rect 1082 -924 1088 -864
rect 2052 -924 2058 -864
rect 2118 -924 2124 -864
rect 2186 -1034 2246 -804
rect 2314 -1034 2374 -804
rect 656 -1066 2434 -1034
rect 656 -1134 692 -1066
rect 2400 -1134 2434 -1066
rect 656 -1164 2434 -1134
rect 432 -1616 544 -1530
rect 1144 -1616 1154 -1316
rect 2046 -1616 2056 -1316
rect 2656 -1530 2662 130
rect 2762 -1530 2768 130
rect 2656 -1616 2768 -1530
rect 432 -1622 2768 -1616
rect 432 -1722 538 -1622
rect 2662 -1722 2768 -1622
rect 432 -1728 2768 -1722
<< via1 >>
rect 544 3256 1144 3556
rect 2056 3256 2656 3556
rect 734 2988 2558 3052
rect 1288 2814 1348 2874
rect 1806 2814 1866 2874
rect 626 2582 686 2642
rect 626 1988 686 2048
rect 1160 1858 1220 1918
rect 1030 1744 1090 1804
rect 876 1008 936 1068
rect 1544 2702 1604 2762
rect 1416 2582 1476 2642
rect 1672 2582 1732 2642
rect 2474 2702 2534 2762
rect 1418 1858 1478 1918
rect 1676 1858 1736 1918
rect 1548 1744 1608 1804
rect 1934 1858 1994 1918
rect 2064 1744 2124 1804
rect 1160 1008 1220 1068
rect 1028 896 1088 956
rect 1936 1008 1996 1068
rect 2064 896 2124 956
rect 1544 748 1604 808
rect 1802 788 1862 848
rect 2474 896 2534 956
rect -108 472 -48 532
rect 214 468 274 474
rect 214 420 220 468
rect 220 420 268 468
rect 268 420 274 468
rect 214 414 274 420
rect 1544 108 1604 168
rect 1028 42 1088 102
rect 1282 -2 1342 58
rect 1414 -114 1474 -54
rect 1802 -2 1862 58
rect 1670 -114 1730 -54
rect 1156 -810 1216 -750
rect 1930 -810 1990 -750
rect 1022 -924 1082 -864
rect 2058 -924 2118 -864
rect 692 -1134 2400 -1066
rect 544 -1616 1144 -1316
rect 2056 -1616 2656 -1316
<< metal2 >>
rect 544 3556 1144 3566
rect 544 3246 1144 3256
rect 2056 3556 2656 3566
rect 2056 3246 2656 3256
rect 700 3052 2602 3082
rect 700 2988 734 3052
rect 2558 2988 2602 3052
rect 700 2958 2602 2988
rect 1288 2874 1348 2880
rect 1806 2874 1866 2880
rect 1348 2814 1806 2874
rect 1288 2808 1348 2814
rect 1806 2808 1866 2814
rect 1544 2762 1604 2768
rect 2474 2762 2534 2768
rect 1604 2702 2474 2762
rect 1544 2696 1604 2702
rect 2474 2696 2534 2702
rect 626 2642 686 2648
rect 1416 2642 1476 2648
rect 1672 2642 1732 2648
rect 686 2582 1416 2642
rect 1476 2582 1672 2642
rect 626 2576 686 2582
rect 1416 2576 1476 2582
rect 1672 2576 1732 2582
rect -108 1988 626 2048
rect 686 1988 692 2048
rect -108 532 -48 1988
rect 1160 1918 1220 1924
rect 1418 1918 1478 1924
rect 1676 1918 1736 1924
rect 1934 1918 1994 1924
rect 628 1858 1160 1918
rect 1220 1858 1418 1918
rect 1478 1858 1676 1918
rect 1736 1858 1934 1918
rect -114 472 -108 532
rect -48 472 -42 532
rect 628 474 688 1858
rect 1160 1852 1220 1858
rect 1418 1852 1478 1858
rect 1676 1852 1736 1858
rect 1934 1852 1994 1858
rect 1030 1804 1090 1810
rect 1548 1804 1608 1810
rect 2064 1804 2124 1810
rect 1090 1744 1548 1804
rect 1608 1744 2064 1804
rect 1030 1738 1090 1744
rect 1548 1738 1608 1744
rect 2064 1738 2124 1744
rect 208 414 214 474
rect 274 414 688 474
rect 628 -750 688 414
rect 876 1068 936 1074
rect 1160 1068 1220 1074
rect 1936 1068 1996 1074
rect 936 1008 1160 1068
rect 1220 1008 1936 1068
rect 876 -54 936 1008
rect 1160 1002 1220 1008
rect 1936 1002 1996 1008
rect 1028 956 1088 962
rect 2064 956 2124 962
rect 2474 956 2534 962
rect 1088 896 2064 956
rect 2124 896 2474 956
rect 1028 102 1088 896
rect 2064 890 2124 896
rect 2474 890 2534 896
rect 1802 848 1862 854
rect 1544 808 1604 814
rect 1544 168 1604 748
rect 1538 108 1544 168
rect 1604 108 1610 168
rect 1028 36 1088 42
rect 1282 58 1342 64
rect 1802 58 1862 788
rect 1342 -2 1802 58
rect 1282 -8 1342 -2
rect 1802 -8 1862 -2
rect 1414 -54 1474 -48
rect 1670 -54 1730 -48
rect 876 -114 1414 -54
rect 1474 -114 1670 -54
rect 1414 -120 1474 -114
rect 1670 -120 1730 -114
rect 1156 -750 1216 -744
rect 1930 -750 1990 -744
rect 628 -810 1156 -750
rect 1216 -810 1930 -750
rect 1156 -816 1216 -810
rect 1930 -816 1990 -810
rect 1022 -864 1082 -858
rect 2058 -864 2118 -858
rect 1082 -924 2058 -864
rect 1022 -930 1082 -924
rect 2058 -930 2118 -924
rect 656 -1066 2434 -1034
rect 656 -1134 692 -1066
rect 2400 -1134 2434 -1066
rect 656 -1164 2434 -1134
rect 544 -1316 1144 -1306
rect 544 -1626 1144 -1616
rect 2056 -1316 2656 -1306
rect 2056 -1626 2656 -1616
<< via2 >>
rect 544 3256 1144 3556
rect 2056 3256 2656 3556
rect 734 2988 2558 3052
rect 692 -1134 2400 -1066
rect 544 -1616 1144 -1316
rect 2056 -1616 2656 -1316
<< metal3 >>
rect 534 3556 1154 3561
rect 534 3256 544 3556
rect 1144 3256 1154 3556
rect 534 3251 1154 3256
rect 2046 3556 2666 3561
rect 2046 3256 2056 3556
rect 2656 3256 2666 3556
rect 2046 3251 2666 3256
rect 700 3052 2602 3082
rect 700 2988 734 3052
rect 2558 2988 2602 3052
rect 700 2958 2602 2988
rect 656 -1066 2434 -1034
rect 656 -1134 692 -1066
rect 2400 -1134 2434 -1066
rect 656 -1164 2434 -1134
rect 534 -1316 1154 -1311
rect 534 -1616 544 -1316
rect 1144 -1616 1154 -1316
rect 534 -1621 1154 -1616
rect 2046 -1316 2666 -1311
rect 2046 -1616 2056 -1316
rect 2656 -1616 2666 -1316
rect 2046 -1621 2666 -1616
<< via3 >>
rect 544 3256 1144 3556
rect 2056 3256 2656 3556
rect 734 2988 2558 3052
rect 692 -1134 2400 -1066
rect 544 -1616 1144 -1316
rect 2056 -1616 2656 -1316
<< metal4 >>
rect 360 3556 2840 3740
rect 360 3256 544 3556
rect 1144 3256 2056 3556
rect 2656 3256 2840 3556
rect 360 3052 2840 3256
rect 360 2988 734 3052
rect 2558 2988 2840 3052
rect 360 2940 2840 2988
rect 360 -1066 2840 -1000
rect 360 -1134 692 -1066
rect 2400 -1134 2840 -1066
rect 360 -1316 2840 -1134
rect 360 -1616 544 -1316
rect 1144 -1616 2056 -1316
rect 2656 -1616 2840 -1316
rect 360 -1800 2840 -1616
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623971255
transform 1 0 50 0 1 262
box -38 -48 314 592
use sky130_fd_pr__nfet_01v8_V7QVDJ  sky130_fd_pr__nfet_01v8_V7QVDJ_0
timestamp 1623971255
transform 1 0 1571 0 1 -430
box -803 -288 803 288
use sky130_fd_pr__pfet_01v8_hvt_RC2PSP  sky130_fd_pr__pfet_01v8_hvt_RC2PSP_1
timestamp 1623971255
transform 1 0 1576 0 1 2263
box -839 -300 839 300
use sky130_fd_pr__pfet_01v8_hvt_RC2PSP  sky130_fd_pr__pfet_01v8_hvt_RC2PSP_0
timestamp 1623971255
transform 1 0 1576 0 1 1403
box -839 -300 839 300
<< labels >>
flabel metal1 -26 494 -20 498 1 FreeSans 480 0 0 0 SEL
flabel metal2 1570 420 1578 428 1 FreeSans 480 0 0 0 A
flabel metal2 1824 440 1832 446 1 FreeSans 480 0 0 0 Y
flabel metal2 1048 442 1058 448 1 FreeSans 480 0 0 0 B
flabel metal2 434 442 444 452 1 FreeSans 480 0 0 0 SELB
flabel metal4 1310 3714 1322 3724 1 FreeSans 480 0 0 0 VDD
flabel metal4 1382 -1784 1396 -1776 1 FreeSans 480 0 0 0 VSS
<< properties >>
string FIXED_BBOX 488 -1672 2712 272
<< end >>

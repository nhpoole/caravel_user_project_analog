magic
tech sky130A
magscale 1 2
timestamp 1624298412
<< nwell >>
rect 342 -10384 24858 4358
<< pwell >>
rect -12358 -27258 24958 -11142
<< nmos >>
rect 2628 -14832 3588 -14232
rect 3646 -14832 4606 -14232
rect 4664 -14832 5624 -14232
rect 5682 -14832 6642 -14232
rect 6700 -14832 7660 -14232
rect 7718 -14832 8678 -14232
rect 8736 -14832 9696 -14232
rect 9754 -14832 10714 -14232
rect 10772 -14832 11732 -14232
rect 11790 -14832 12750 -14232
rect 12808 -14832 13768 -14232
rect 13826 -14832 14786 -14232
rect 14844 -14832 15804 -14232
rect 15862 -14832 16822 -14232
rect 16880 -14832 17840 -14232
rect 17898 -14832 18858 -14232
rect 18916 -14832 19876 -14232
rect 19934 -14832 20894 -14232
rect 20952 -14832 21912 -14232
rect 21970 -14832 22930 -14232
rect 2628 -16064 3588 -15464
rect 3646 -16064 4606 -15464
rect 4664 -16064 5624 -15464
rect 5682 -16064 6642 -15464
rect 6700 -16064 7660 -15464
rect 7718 -16064 8678 -15464
rect 8736 -16064 9696 -15464
rect 9754 -16064 10714 -15464
rect 10772 -16064 11732 -15464
rect 11790 -16064 12750 -15464
rect 12808 -16064 13768 -15464
rect 13826 -16064 14786 -15464
rect 14844 -16064 15804 -15464
rect 15862 -16064 16822 -15464
rect 16880 -16064 17840 -15464
rect 17898 -16064 18858 -15464
rect 18916 -16064 19876 -15464
rect 19934 -16064 20894 -15464
rect 20952 -16064 21912 -15464
rect 21970 -16064 22930 -15464
rect 2626 -17298 3586 -16698
rect 3644 -17298 4604 -16698
rect 4662 -17298 5622 -16698
rect 5680 -17298 6640 -16698
rect 6698 -17298 7658 -16698
rect 7716 -17298 8676 -16698
rect 8734 -17298 9694 -16698
rect 9752 -17298 10712 -16698
rect 10770 -17298 11730 -16698
rect 11788 -17298 12748 -16698
rect 12806 -17298 13766 -16698
rect 13824 -17298 14784 -16698
rect 14842 -17298 15802 -16698
rect 15860 -17298 16820 -16698
rect 16878 -17298 17838 -16698
rect 17896 -17298 18856 -16698
rect 18914 -17298 19874 -16698
rect 19932 -17298 20892 -16698
rect 20950 -17298 21910 -16698
rect 21968 -17298 22928 -16698
rect 2626 -18532 3586 -17932
rect 3644 -18532 4604 -17932
rect 4662 -18532 5622 -17932
rect 5680 -18532 6640 -17932
rect 6698 -18532 7658 -17932
rect 7716 -18532 8676 -17932
rect 8734 -18532 9694 -17932
rect 9752 -18532 10712 -17932
rect 10770 -18532 11730 -17932
rect 11788 -18532 12748 -17932
rect 12806 -18532 13766 -17932
rect 13824 -18532 14784 -17932
rect 14842 -18532 15802 -17932
rect 15860 -18532 16820 -17932
rect 16878 -18532 17838 -17932
rect 17896 -18532 18856 -17932
rect 18914 -18532 19874 -17932
rect 19932 -18532 20892 -17932
rect 20950 -18532 21910 -17932
rect 21968 -18532 22928 -17932
rect 2626 -19764 3586 -19164
rect 3644 -19764 4604 -19164
rect 4662 -19764 5622 -19164
rect 5680 -19764 6640 -19164
rect 6698 -19764 7658 -19164
rect 7716 -19764 8676 -19164
rect 8734 -19764 9694 -19164
rect 9752 -19764 10712 -19164
rect 10770 -19764 11730 -19164
rect 11788 -19764 12748 -19164
rect 12806 -19764 13766 -19164
rect 13824 -19764 14784 -19164
rect 14842 -19764 15802 -19164
rect 15860 -19764 16820 -19164
rect 16878 -19764 17838 -19164
rect 17896 -19764 18856 -19164
rect 18914 -19764 19874 -19164
rect 19932 -19764 20892 -19164
rect 20950 -19764 21910 -19164
rect 21968 -19764 22928 -19164
rect 2626 -20998 3586 -20398
rect 3644 -20998 4604 -20398
rect 4662 -20998 5622 -20398
rect 5680 -20998 6640 -20398
rect 6698 -20998 7658 -20398
rect 7716 -20998 8676 -20398
rect 8734 -20998 9694 -20398
rect 9752 -20998 10712 -20398
rect 10770 -20998 11730 -20398
rect 11788 -20998 12748 -20398
rect 12806 -20998 13766 -20398
rect 13824 -20998 14784 -20398
rect 14842 -20998 15802 -20398
rect 15860 -20998 16820 -20398
rect 16878 -20998 17838 -20398
rect 17896 -20998 18856 -20398
rect 18914 -20998 19874 -20398
rect 19932 -20998 20892 -20398
rect 20950 -20998 21910 -20398
rect 21968 -20998 22928 -20398
rect 2626 -22232 3586 -21632
rect 3644 -22232 4604 -21632
rect 4662 -22232 5622 -21632
rect 5680 -22232 6640 -21632
rect 6698 -22232 7658 -21632
rect 7716 -22232 8676 -21632
rect 8734 -22232 9694 -21632
rect 9752 -22232 10712 -21632
rect 10770 -22232 11730 -21632
rect 11788 -22232 12748 -21632
rect 12806 -22232 13766 -21632
rect 13824 -22232 14784 -21632
rect 14842 -22232 15802 -21632
rect 15860 -22232 16820 -21632
rect 16878 -22232 17838 -21632
rect 17896 -22232 18856 -21632
rect 18914 -22232 19874 -21632
rect 19932 -22232 20892 -21632
rect 20950 -22232 21910 -21632
rect 21968 -22232 22928 -21632
rect 2626 -23464 3586 -22864
rect 3644 -23464 4604 -22864
rect 4662 -23464 5622 -22864
rect 5680 -23464 6640 -22864
rect 6698 -23464 7658 -22864
rect 7716 -23464 8676 -22864
rect 8734 -23464 9694 -22864
rect 9752 -23464 10712 -22864
rect 10770 -23464 11730 -22864
rect 11788 -23464 12748 -22864
rect 12806 -23464 13766 -22864
rect 13824 -23464 14784 -22864
rect 14842 -23464 15802 -22864
rect 15860 -23464 16820 -22864
rect 16878 -23464 17838 -22864
rect 17896 -23464 18856 -22864
rect 18914 -23464 19874 -22864
rect 19932 -23464 20892 -22864
rect 20950 -23464 21910 -22864
rect 21968 -23464 22928 -22864
rect 2626 -24698 3586 -24098
rect 3644 -24698 4604 -24098
rect 4662 -24698 5622 -24098
rect 5680 -24698 6640 -24098
rect 6698 -24698 7658 -24098
rect 7716 -24698 8676 -24098
rect 8734 -24698 9694 -24098
rect 9752 -24698 10712 -24098
rect 10770 -24698 11730 -24098
rect 11788 -24698 12748 -24098
rect 12806 -24698 13766 -24098
rect 13824 -24698 14784 -24098
rect 14842 -24698 15802 -24098
rect 15860 -24698 16820 -24098
rect 16878 -24698 17838 -24098
rect 17896 -24698 18856 -24098
rect 18914 -24698 19874 -24098
rect 19932 -24698 20892 -24098
rect 20950 -24698 21910 -24098
rect 21968 -24698 22928 -24098
<< nmoslvt >>
rect -9138 -13112 -8178 -12512
rect -8120 -13112 -7160 -12512
rect -7102 -13112 -6142 -12512
rect -6084 -13112 -5124 -12512
rect -5066 -13112 -4106 -12512
rect -4048 -13112 -3088 -12512
rect -3030 -13112 -2070 -12512
rect -2012 -13112 -1052 -12512
rect -994 -13112 -34 -12512
rect -9138 -13930 -8178 -13330
rect -8120 -13930 -7160 -13330
rect -7102 -13930 -6142 -13330
rect -6084 -13930 -5124 -13330
rect -5066 -13930 -4106 -13330
rect -4048 -13930 -3088 -13330
rect -3030 -13930 -2070 -13330
rect -2012 -13930 -1052 -13330
rect -994 -13930 -34 -13330
rect -9138 -14748 -8178 -14148
rect -8120 -14748 -7160 -14148
rect -7102 -14748 -6142 -14148
rect -6084 -14748 -5124 -14148
rect -5066 -14748 -4106 -14148
rect -4048 -14748 -3088 -14148
rect -3030 -14748 -2070 -14148
rect -2012 -14748 -1052 -14148
rect -994 -14748 -34 -14148
rect -9138 -15566 -8178 -14966
rect -8120 -15566 -7160 -14966
rect -7102 -15566 -6142 -14966
rect -6084 -15566 -5124 -14966
rect -5066 -15566 -4106 -14966
rect -4048 -15566 -3088 -14966
rect -3030 -15566 -2070 -14966
rect -2012 -15566 -1052 -14966
rect -994 -15566 -34 -14966
rect -9138 -16384 -8178 -15784
rect -8120 -16384 -7160 -15784
rect -7102 -16384 -6142 -15784
rect -6084 -16384 -5124 -15784
rect -5066 -16384 -4106 -15784
rect -4048 -16384 -3088 -15784
rect -3030 -16384 -2070 -15784
rect -2012 -16384 -1052 -15784
rect -994 -16384 -34 -15784
rect -9138 -17202 -8178 -16602
rect -8120 -17202 -7160 -16602
rect -7102 -17202 -6142 -16602
rect -6084 -17202 -5124 -16602
rect -5066 -17202 -4106 -16602
rect -4048 -17202 -3088 -16602
rect -3030 -17202 -2070 -16602
rect -2012 -17202 -1052 -16602
rect -994 -17202 -34 -16602
rect -9138 -18020 -8178 -17420
rect -8120 -18020 -7160 -17420
rect -7102 -18020 -6142 -17420
rect -6084 -18020 -5124 -17420
rect -5066 -18020 -4106 -17420
rect -4048 -18020 -3088 -17420
rect -3030 -18020 -2070 -17420
rect -2012 -18020 -1052 -17420
rect -994 -18020 -34 -17420
rect -9138 -18838 -8178 -18238
rect -8120 -18838 -7160 -18238
rect -7102 -18838 -6142 -18238
rect -6084 -18838 -5124 -18238
rect -5066 -18838 -4106 -18238
rect -4048 -18838 -3088 -18238
rect -3030 -18838 -2070 -18238
rect -2012 -18838 -1052 -18238
rect -994 -18838 -34 -18238
<< ndiff >>
rect -9196 -12524 -9138 -12512
rect -9196 -13100 -9184 -12524
rect -9150 -13100 -9138 -12524
rect -9196 -13112 -9138 -13100
rect -8178 -12524 -8120 -12512
rect -8178 -13100 -8166 -12524
rect -8132 -13100 -8120 -12524
rect -8178 -13112 -8120 -13100
rect -7160 -12524 -7102 -12512
rect -7160 -13100 -7148 -12524
rect -7114 -13100 -7102 -12524
rect -7160 -13112 -7102 -13100
rect -6142 -12524 -6084 -12512
rect -6142 -13100 -6130 -12524
rect -6096 -13100 -6084 -12524
rect -6142 -13112 -6084 -13100
rect -5124 -12524 -5066 -12512
rect -5124 -13100 -5112 -12524
rect -5078 -13100 -5066 -12524
rect -5124 -13112 -5066 -13100
rect -4106 -12524 -4048 -12512
rect -4106 -13100 -4094 -12524
rect -4060 -13100 -4048 -12524
rect -4106 -13112 -4048 -13100
rect -3088 -12524 -3030 -12512
rect -3088 -13100 -3076 -12524
rect -3042 -13100 -3030 -12524
rect -3088 -13112 -3030 -13100
rect -2070 -12524 -2012 -12512
rect -2070 -13100 -2058 -12524
rect -2024 -13100 -2012 -12524
rect -2070 -13112 -2012 -13100
rect -1052 -12524 -994 -12512
rect -1052 -13100 -1040 -12524
rect -1006 -13100 -994 -12524
rect -1052 -13112 -994 -13100
rect -34 -12524 24 -12512
rect -34 -13100 -22 -12524
rect 12 -13100 24 -12524
rect -34 -13112 24 -13100
rect -9196 -13342 -9138 -13330
rect -9196 -13918 -9184 -13342
rect -9150 -13918 -9138 -13342
rect -9196 -13930 -9138 -13918
rect -8178 -13342 -8120 -13330
rect -8178 -13918 -8166 -13342
rect -8132 -13918 -8120 -13342
rect -8178 -13930 -8120 -13918
rect -7160 -13342 -7102 -13330
rect -7160 -13918 -7148 -13342
rect -7114 -13918 -7102 -13342
rect -7160 -13930 -7102 -13918
rect -6142 -13342 -6084 -13330
rect -6142 -13918 -6130 -13342
rect -6096 -13918 -6084 -13342
rect -6142 -13930 -6084 -13918
rect -5124 -13342 -5066 -13330
rect -5124 -13918 -5112 -13342
rect -5078 -13918 -5066 -13342
rect -5124 -13930 -5066 -13918
rect -4106 -13342 -4048 -13330
rect -4106 -13918 -4094 -13342
rect -4060 -13918 -4048 -13342
rect -4106 -13930 -4048 -13918
rect -3088 -13342 -3030 -13330
rect -3088 -13918 -3076 -13342
rect -3042 -13918 -3030 -13342
rect -3088 -13930 -3030 -13918
rect -2070 -13342 -2012 -13330
rect -2070 -13918 -2058 -13342
rect -2024 -13918 -2012 -13342
rect -2070 -13930 -2012 -13918
rect -1052 -13342 -994 -13330
rect -1052 -13918 -1040 -13342
rect -1006 -13918 -994 -13342
rect -1052 -13930 -994 -13918
rect -34 -13342 24 -13330
rect -34 -13918 -22 -13342
rect 12 -13918 24 -13342
rect -34 -13930 24 -13918
rect -9196 -14160 -9138 -14148
rect -9196 -14736 -9184 -14160
rect -9150 -14736 -9138 -14160
rect -9196 -14748 -9138 -14736
rect -8178 -14160 -8120 -14148
rect -8178 -14736 -8166 -14160
rect -8132 -14736 -8120 -14160
rect -8178 -14748 -8120 -14736
rect -7160 -14160 -7102 -14148
rect -7160 -14736 -7148 -14160
rect -7114 -14736 -7102 -14160
rect -7160 -14748 -7102 -14736
rect -6142 -14160 -6084 -14148
rect -6142 -14736 -6130 -14160
rect -6096 -14736 -6084 -14160
rect -6142 -14748 -6084 -14736
rect -5124 -14160 -5066 -14148
rect -5124 -14736 -5112 -14160
rect -5078 -14736 -5066 -14160
rect -5124 -14748 -5066 -14736
rect -4106 -14160 -4048 -14148
rect -4106 -14736 -4094 -14160
rect -4060 -14736 -4048 -14160
rect -4106 -14748 -4048 -14736
rect -3088 -14160 -3030 -14148
rect -3088 -14736 -3076 -14160
rect -3042 -14736 -3030 -14160
rect -3088 -14748 -3030 -14736
rect -2070 -14160 -2012 -14148
rect -2070 -14736 -2058 -14160
rect -2024 -14736 -2012 -14160
rect -2070 -14748 -2012 -14736
rect -1052 -14160 -994 -14148
rect -1052 -14736 -1040 -14160
rect -1006 -14736 -994 -14160
rect -1052 -14748 -994 -14736
rect -34 -14160 24 -14148
rect -34 -14736 -22 -14160
rect 12 -14736 24 -14160
rect -34 -14748 24 -14736
rect 2570 -14244 2628 -14232
rect 2570 -14820 2582 -14244
rect 2616 -14820 2628 -14244
rect 2570 -14832 2628 -14820
rect 3588 -14244 3646 -14232
rect 3588 -14820 3600 -14244
rect 3634 -14820 3646 -14244
rect 3588 -14832 3646 -14820
rect 4606 -14244 4664 -14232
rect 4606 -14820 4618 -14244
rect 4652 -14820 4664 -14244
rect 4606 -14832 4664 -14820
rect 5624 -14244 5682 -14232
rect 5624 -14820 5636 -14244
rect 5670 -14820 5682 -14244
rect 5624 -14832 5682 -14820
rect 6642 -14244 6700 -14232
rect 6642 -14820 6654 -14244
rect 6688 -14820 6700 -14244
rect 6642 -14832 6700 -14820
rect 7660 -14244 7718 -14232
rect 7660 -14820 7672 -14244
rect 7706 -14820 7718 -14244
rect 7660 -14832 7718 -14820
rect 8678 -14244 8736 -14232
rect 8678 -14820 8690 -14244
rect 8724 -14820 8736 -14244
rect 8678 -14832 8736 -14820
rect 9696 -14244 9754 -14232
rect 9696 -14820 9708 -14244
rect 9742 -14820 9754 -14244
rect 9696 -14832 9754 -14820
rect 10714 -14244 10772 -14232
rect 10714 -14820 10726 -14244
rect 10760 -14820 10772 -14244
rect 10714 -14832 10772 -14820
rect 11732 -14244 11790 -14232
rect 11732 -14820 11744 -14244
rect 11778 -14820 11790 -14244
rect 11732 -14832 11790 -14820
rect 12750 -14244 12808 -14232
rect 12750 -14820 12762 -14244
rect 12796 -14820 12808 -14244
rect 12750 -14832 12808 -14820
rect 13768 -14244 13826 -14232
rect 13768 -14820 13780 -14244
rect 13814 -14820 13826 -14244
rect 13768 -14832 13826 -14820
rect 14786 -14244 14844 -14232
rect 14786 -14820 14798 -14244
rect 14832 -14820 14844 -14244
rect 14786 -14832 14844 -14820
rect 15804 -14244 15862 -14232
rect 15804 -14820 15816 -14244
rect 15850 -14820 15862 -14244
rect 15804 -14832 15862 -14820
rect 16822 -14244 16880 -14232
rect 16822 -14820 16834 -14244
rect 16868 -14820 16880 -14244
rect 16822 -14832 16880 -14820
rect 17840 -14244 17898 -14232
rect 17840 -14820 17852 -14244
rect 17886 -14820 17898 -14244
rect 17840 -14832 17898 -14820
rect 18858 -14244 18916 -14232
rect 18858 -14820 18870 -14244
rect 18904 -14820 18916 -14244
rect 18858 -14832 18916 -14820
rect 19876 -14244 19934 -14232
rect 19876 -14820 19888 -14244
rect 19922 -14820 19934 -14244
rect 19876 -14832 19934 -14820
rect 20894 -14244 20952 -14232
rect 20894 -14820 20906 -14244
rect 20940 -14820 20952 -14244
rect 20894 -14832 20952 -14820
rect 21912 -14244 21970 -14232
rect 21912 -14820 21924 -14244
rect 21958 -14820 21970 -14244
rect 21912 -14832 21970 -14820
rect 22930 -14244 22988 -14232
rect 22930 -14820 22942 -14244
rect 22976 -14820 22988 -14244
rect 22930 -14832 22988 -14820
rect -9196 -14978 -9138 -14966
rect -9196 -15554 -9184 -14978
rect -9150 -15554 -9138 -14978
rect -9196 -15566 -9138 -15554
rect -8178 -14978 -8120 -14966
rect -8178 -15554 -8166 -14978
rect -8132 -15554 -8120 -14978
rect -8178 -15566 -8120 -15554
rect -7160 -14978 -7102 -14966
rect -7160 -15554 -7148 -14978
rect -7114 -15554 -7102 -14978
rect -7160 -15566 -7102 -15554
rect -6142 -14978 -6084 -14966
rect -6142 -15554 -6130 -14978
rect -6096 -15554 -6084 -14978
rect -6142 -15566 -6084 -15554
rect -5124 -14978 -5066 -14966
rect -5124 -15554 -5112 -14978
rect -5078 -15554 -5066 -14978
rect -5124 -15566 -5066 -15554
rect -4106 -14978 -4048 -14966
rect -4106 -15554 -4094 -14978
rect -4060 -15554 -4048 -14978
rect -4106 -15566 -4048 -15554
rect -3088 -14978 -3030 -14966
rect -3088 -15554 -3076 -14978
rect -3042 -15554 -3030 -14978
rect -3088 -15566 -3030 -15554
rect -2070 -14978 -2012 -14966
rect -2070 -15554 -2058 -14978
rect -2024 -15554 -2012 -14978
rect -2070 -15566 -2012 -15554
rect -1052 -14978 -994 -14966
rect -1052 -15554 -1040 -14978
rect -1006 -15554 -994 -14978
rect -1052 -15566 -994 -15554
rect -34 -14978 24 -14966
rect -34 -15554 -22 -14978
rect 12 -15554 24 -14978
rect -34 -15566 24 -15554
rect 2570 -15476 2628 -15464
rect -9196 -15796 -9138 -15784
rect -9196 -16372 -9184 -15796
rect -9150 -16372 -9138 -15796
rect -9196 -16384 -9138 -16372
rect -8178 -15796 -8120 -15784
rect -8178 -16372 -8166 -15796
rect -8132 -16372 -8120 -15796
rect -8178 -16384 -8120 -16372
rect -7160 -15796 -7102 -15784
rect -7160 -16372 -7148 -15796
rect -7114 -16372 -7102 -15796
rect -7160 -16384 -7102 -16372
rect -6142 -15796 -6084 -15784
rect -6142 -16372 -6130 -15796
rect -6096 -16372 -6084 -15796
rect -6142 -16384 -6084 -16372
rect -5124 -15796 -5066 -15784
rect -5124 -16372 -5112 -15796
rect -5078 -16372 -5066 -15796
rect -5124 -16384 -5066 -16372
rect -4106 -15796 -4048 -15784
rect -4106 -16372 -4094 -15796
rect -4060 -16372 -4048 -15796
rect -4106 -16384 -4048 -16372
rect -3088 -15796 -3030 -15784
rect -3088 -16372 -3076 -15796
rect -3042 -16372 -3030 -15796
rect -3088 -16384 -3030 -16372
rect -2070 -15796 -2012 -15784
rect -2070 -16372 -2058 -15796
rect -2024 -16372 -2012 -15796
rect -2070 -16384 -2012 -16372
rect -1052 -15796 -994 -15784
rect -1052 -16372 -1040 -15796
rect -1006 -16372 -994 -15796
rect -1052 -16384 -994 -16372
rect -34 -15796 24 -15784
rect -34 -16372 -22 -15796
rect 12 -16372 24 -15796
rect 2570 -16052 2582 -15476
rect 2616 -16052 2628 -15476
rect 2570 -16064 2628 -16052
rect 3588 -15476 3646 -15464
rect 3588 -16052 3600 -15476
rect 3634 -16052 3646 -15476
rect 3588 -16064 3646 -16052
rect 4606 -15476 4664 -15464
rect 4606 -16052 4618 -15476
rect 4652 -16052 4664 -15476
rect 4606 -16064 4664 -16052
rect 5624 -15476 5682 -15464
rect 5624 -16052 5636 -15476
rect 5670 -16052 5682 -15476
rect 5624 -16064 5682 -16052
rect 6642 -15476 6700 -15464
rect 6642 -16052 6654 -15476
rect 6688 -16052 6700 -15476
rect 6642 -16064 6700 -16052
rect 7660 -15476 7718 -15464
rect 7660 -16052 7672 -15476
rect 7706 -16052 7718 -15476
rect 7660 -16064 7718 -16052
rect 8678 -15476 8736 -15464
rect 8678 -16052 8690 -15476
rect 8724 -16052 8736 -15476
rect 8678 -16064 8736 -16052
rect 9696 -15476 9754 -15464
rect 9696 -16052 9708 -15476
rect 9742 -16052 9754 -15476
rect 9696 -16064 9754 -16052
rect 10714 -15476 10772 -15464
rect 10714 -16052 10726 -15476
rect 10760 -16052 10772 -15476
rect 10714 -16064 10772 -16052
rect 11732 -15476 11790 -15464
rect 11732 -16052 11744 -15476
rect 11778 -16052 11790 -15476
rect 11732 -16064 11790 -16052
rect 12750 -15476 12808 -15464
rect 12750 -16052 12762 -15476
rect 12796 -16052 12808 -15476
rect 12750 -16064 12808 -16052
rect 13768 -15476 13826 -15464
rect 13768 -16052 13780 -15476
rect 13814 -16052 13826 -15476
rect 13768 -16064 13826 -16052
rect 14786 -15476 14844 -15464
rect 14786 -16052 14798 -15476
rect 14832 -16052 14844 -15476
rect 14786 -16064 14844 -16052
rect 15804 -15476 15862 -15464
rect 15804 -16052 15816 -15476
rect 15850 -16052 15862 -15476
rect 15804 -16064 15862 -16052
rect 16822 -15476 16880 -15464
rect 16822 -16052 16834 -15476
rect 16868 -16052 16880 -15476
rect 16822 -16064 16880 -16052
rect 17840 -15476 17898 -15464
rect 17840 -16052 17852 -15476
rect 17886 -16052 17898 -15476
rect 17840 -16064 17898 -16052
rect 18858 -15476 18916 -15464
rect 18858 -16052 18870 -15476
rect 18904 -16052 18916 -15476
rect 18858 -16064 18916 -16052
rect 19876 -15476 19934 -15464
rect 19876 -16052 19888 -15476
rect 19922 -16052 19934 -15476
rect 19876 -16064 19934 -16052
rect 20894 -15476 20952 -15464
rect 20894 -16052 20906 -15476
rect 20940 -16052 20952 -15476
rect 20894 -16064 20952 -16052
rect 21912 -15476 21970 -15464
rect 21912 -16052 21924 -15476
rect 21958 -16052 21970 -15476
rect 21912 -16064 21970 -16052
rect 22930 -15476 22988 -15464
rect 22930 -16052 22942 -15476
rect 22976 -16052 22988 -15476
rect 22930 -16064 22988 -16052
rect -34 -16384 24 -16372
rect -9196 -16614 -9138 -16602
rect -9196 -17190 -9184 -16614
rect -9150 -17190 -9138 -16614
rect -9196 -17202 -9138 -17190
rect -8178 -16614 -8120 -16602
rect -8178 -17190 -8166 -16614
rect -8132 -17190 -8120 -16614
rect -8178 -17202 -8120 -17190
rect -7160 -16614 -7102 -16602
rect -7160 -17190 -7148 -16614
rect -7114 -17190 -7102 -16614
rect -7160 -17202 -7102 -17190
rect -6142 -16614 -6084 -16602
rect -6142 -17190 -6130 -16614
rect -6096 -17190 -6084 -16614
rect -6142 -17202 -6084 -17190
rect -5124 -16614 -5066 -16602
rect -5124 -17190 -5112 -16614
rect -5078 -17190 -5066 -16614
rect -5124 -17202 -5066 -17190
rect -4106 -16614 -4048 -16602
rect -4106 -17190 -4094 -16614
rect -4060 -17190 -4048 -16614
rect -4106 -17202 -4048 -17190
rect -3088 -16614 -3030 -16602
rect -3088 -17190 -3076 -16614
rect -3042 -17190 -3030 -16614
rect -3088 -17202 -3030 -17190
rect -2070 -16614 -2012 -16602
rect -2070 -17190 -2058 -16614
rect -2024 -17190 -2012 -16614
rect -2070 -17202 -2012 -17190
rect -1052 -16614 -994 -16602
rect -1052 -17190 -1040 -16614
rect -1006 -17190 -994 -16614
rect -1052 -17202 -994 -17190
rect -34 -16614 24 -16602
rect -34 -17190 -22 -16614
rect 12 -17190 24 -16614
rect -34 -17202 24 -17190
rect 2568 -16710 2626 -16698
rect 2568 -17286 2580 -16710
rect 2614 -17286 2626 -16710
rect 2568 -17298 2626 -17286
rect 3586 -16710 3644 -16698
rect 3586 -17286 3598 -16710
rect 3632 -17286 3644 -16710
rect 3586 -17298 3644 -17286
rect 4604 -16710 4662 -16698
rect 4604 -17286 4616 -16710
rect 4650 -17286 4662 -16710
rect 4604 -17298 4662 -17286
rect 5622 -16710 5680 -16698
rect 5622 -17286 5634 -16710
rect 5668 -17286 5680 -16710
rect 5622 -17298 5680 -17286
rect 6640 -16710 6698 -16698
rect 6640 -17286 6652 -16710
rect 6686 -17286 6698 -16710
rect 6640 -17298 6698 -17286
rect 7658 -16710 7716 -16698
rect 7658 -17286 7670 -16710
rect 7704 -17286 7716 -16710
rect 7658 -17298 7716 -17286
rect 8676 -16710 8734 -16698
rect 8676 -17286 8688 -16710
rect 8722 -17286 8734 -16710
rect 8676 -17298 8734 -17286
rect 9694 -16710 9752 -16698
rect 9694 -17286 9706 -16710
rect 9740 -17286 9752 -16710
rect 9694 -17298 9752 -17286
rect 10712 -16710 10770 -16698
rect 10712 -17286 10724 -16710
rect 10758 -17286 10770 -16710
rect 10712 -17298 10770 -17286
rect 11730 -16710 11788 -16698
rect 11730 -17286 11742 -16710
rect 11776 -17286 11788 -16710
rect 11730 -17298 11788 -17286
rect 12748 -16710 12806 -16698
rect 12748 -17286 12760 -16710
rect 12794 -17286 12806 -16710
rect 12748 -17298 12806 -17286
rect 13766 -16710 13824 -16698
rect 13766 -17286 13778 -16710
rect 13812 -17286 13824 -16710
rect 13766 -17298 13824 -17286
rect 14784 -16710 14842 -16698
rect 14784 -17286 14796 -16710
rect 14830 -17286 14842 -16710
rect 14784 -17298 14842 -17286
rect 15802 -16710 15860 -16698
rect 15802 -17286 15814 -16710
rect 15848 -17286 15860 -16710
rect 15802 -17298 15860 -17286
rect 16820 -16710 16878 -16698
rect 16820 -17286 16832 -16710
rect 16866 -17286 16878 -16710
rect 16820 -17298 16878 -17286
rect 17838 -16710 17896 -16698
rect 17838 -17286 17850 -16710
rect 17884 -17286 17896 -16710
rect 17838 -17298 17896 -17286
rect 18856 -16710 18914 -16698
rect 18856 -17286 18868 -16710
rect 18902 -17286 18914 -16710
rect 18856 -17298 18914 -17286
rect 19874 -16710 19932 -16698
rect 19874 -17286 19886 -16710
rect 19920 -17286 19932 -16710
rect 19874 -17298 19932 -17286
rect 20892 -16710 20950 -16698
rect 20892 -17286 20904 -16710
rect 20938 -17286 20950 -16710
rect 20892 -17298 20950 -17286
rect 21910 -16710 21968 -16698
rect 21910 -17286 21922 -16710
rect 21956 -17286 21968 -16710
rect 21910 -17298 21968 -17286
rect 22928 -16710 22986 -16698
rect 22928 -17286 22940 -16710
rect 22974 -17286 22986 -16710
rect 22928 -17298 22986 -17286
rect -9196 -17432 -9138 -17420
rect -9196 -18008 -9184 -17432
rect -9150 -18008 -9138 -17432
rect -9196 -18020 -9138 -18008
rect -8178 -17432 -8120 -17420
rect -8178 -18008 -8166 -17432
rect -8132 -18008 -8120 -17432
rect -8178 -18020 -8120 -18008
rect -7160 -17432 -7102 -17420
rect -7160 -18008 -7148 -17432
rect -7114 -18008 -7102 -17432
rect -7160 -18020 -7102 -18008
rect -6142 -17432 -6084 -17420
rect -6142 -18008 -6130 -17432
rect -6096 -18008 -6084 -17432
rect -6142 -18020 -6084 -18008
rect -5124 -17432 -5066 -17420
rect -5124 -18008 -5112 -17432
rect -5078 -18008 -5066 -17432
rect -5124 -18020 -5066 -18008
rect -4106 -17432 -4048 -17420
rect -4106 -18008 -4094 -17432
rect -4060 -18008 -4048 -17432
rect -4106 -18020 -4048 -18008
rect -3088 -17432 -3030 -17420
rect -3088 -18008 -3076 -17432
rect -3042 -18008 -3030 -17432
rect -3088 -18020 -3030 -18008
rect -2070 -17432 -2012 -17420
rect -2070 -18008 -2058 -17432
rect -2024 -18008 -2012 -17432
rect -2070 -18020 -2012 -18008
rect -1052 -17432 -994 -17420
rect -1052 -18008 -1040 -17432
rect -1006 -18008 -994 -17432
rect -1052 -18020 -994 -18008
rect -34 -17432 24 -17420
rect -34 -18008 -22 -17432
rect 12 -18008 24 -17432
rect -34 -18020 24 -18008
rect 2568 -17944 2626 -17932
rect -9196 -18250 -9138 -18238
rect -9196 -18826 -9184 -18250
rect -9150 -18826 -9138 -18250
rect -9196 -18838 -9138 -18826
rect -8178 -18250 -8120 -18238
rect -8178 -18826 -8166 -18250
rect -8132 -18826 -8120 -18250
rect -8178 -18838 -8120 -18826
rect -7160 -18250 -7102 -18238
rect -7160 -18826 -7148 -18250
rect -7114 -18826 -7102 -18250
rect -7160 -18838 -7102 -18826
rect -6142 -18250 -6084 -18238
rect -6142 -18826 -6130 -18250
rect -6096 -18826 -6084 -18250
rect -6142 -18838 -6084 -18826
rect -5124 -18250 -5066 -18238
rect -5124 -18826 -5112 -18250
rect -5078 -18826 -5066 -18250
rect -5124 -18838 -5066 -18826
rect -4106 -18250 -4048 -18238
rect -4106 -18826 -4094 -18250
rect -4060 -18826 -4048 -18250
rect -4106 -18838 -4048 -18826
rect -3088 -18250 -3030 -18238
rect -3088 -18826 -3076 -18250
rect -3042 -18826 -3030 -18250
rect -3088 -18838 -3030 -18826
rect -2070 -18250 -2012 -18238
rect -2070 -18826 -2058 -18250
rect -2024 -18826 -2012 -18250
rect -2070 -18838 -2012 -18826
rect -1052 -18250 -994 -18238
rect -1052 -18826 -1040 -18250
rect -1006 -18826 -994 -18250
rect -1052 -18838 -994 -18826
rect -34 -18250 24 -18238
rect -34 -18826 -22 -18250
rect 12 -18826 24 -18250
rect 2568 -18520 2580 -17944
rect 2614 -18520 2626 -17944
rect 2568 -18532 2626 -18520
rect 3586 -17944 3644 -17932
rect 3586 -18520 3598 -17944
rect 3632 -18520 3644 -17944
rect 3586 -18532 3644 -18520
rect 4604 -17944 4662 -17932
rect 4604 -18520 4616 -17944
rect 4650 -18520 4662 -17944
rect 4604 -18532 4662 -18520
rect 5622 -17944 5680 -17932
rect 5622 -18520 5634 -17944
rect 5668 -18520 5680 -17944
rect 5622 -18532 5680 -18520
rect 6640 -17944 6698 -17932
rect 6640 -18520 6652 -17944
rect 6686 -18520 6698 -17944
rect 6640 -18532 6698 -18520
rect 7658 -17944 7716 -17932
rect 7658 -18520 7670 -17944
rect 7704 -18520 7716 -17944
rect 7658 -18532 7716 -18520
rect 8676 -17944 8734 -17932
rect 8676 -18520 8688 -17944
rect 8722 -18520 8734 -17944
rect 8676 -18532 8734 -18520
rect 9694 -17944 9752 -17932
rect 9694 -18520 9706 -17944
rect 9740 -18520 9752 -17944
rect 9694 -18532 9752 -18520
rect 10712 -17944 10770 -17932
rect 10712 -18520 10724 -17944
rect 10758 -18520 10770 -17944
rect 10712 -18532 10770 -18520
rect 11730 -17944 11788 -17932
rect 11730 -18520 11742 -17944
rect 11776 -18520 11788 -17944
rect 11730 -18532 11788 -18520
rect 12748 -17944 12806 -17932
rect 12748 -18520 12760 -17944
rect 12794 -18520 12806 -17944
rect 12748 -18532 12806 -18520
rect 13766 -17944 13824 -17932
rect 13766 -18520 13778 -17944
rect 13812 -18520 13824 -17944
rect 13766 -18532 13824 -18520
rect 14784 -17944 14842 -17932
rect 14784 -18520 14796 -17944
rect 14830 -18520 14842 -17944
rect 14784 -18532 14842 -18520
rect 15802 -17944 15860 -17932
rect 15802 -18520 15814 -17944
rect 15848 -18520 15860 -17944
rect 15802 -18532 15860 -18520
rect 16820 -17944 16878 -17932
rect 16820 -18520 16832 -17944
rect 16866 -18520 16878 -17944
rect 16820 -18532 16878 -18520
rect 17838 -17944 17896 -17932
rect 17838 -18520 17850 -17944
rect 17884 -18520 17896 -17944
rect 17838 -18532 17896 -18520
rect 18856 -17944 18914 -17932
rect 18856 -18520 18868 -17944
rect 18902 -18520 18914 -17944
rect 18856 -18532 18914 -18520
rect 19874 -17944 19932 -17932
rect 19874 -18520 19886 -17944
rect 19920 -18520 19932 -17944
rect 19874 -18532 19932 -18520
rect 20892 -17944 20950 -17932
rect 20892 -18520 20904 -17944
rect 20938 -18520 20950 -17944
rect 20892 -18532 20950 -18520
rect 21910 -17944 21968 -17932
rect 21910 -18520 21922 -17944
rect 21956 -18520 21968 -17944
rect 21910 -18532 21968 -18520
rect 22928 -17944 22986 -17932
rect 22928 -18520 22940 -17944
rect 22974 -18520 22986 -17944
rect 22928 -18532 22986 -18520
rect -34 -18838 24 -18826
rect 2568 -19176 2626 -19164
rect 2568 -19752 2580 -19176
rect 2614 -19752 2626 -19176
rect 2568 -19764 2626 -19752
rect 3586 -19176 3644 -19164
rect 3586 -19752 3598 -19176
rect 3632 -19752 3644 -19176
rect 3586 -19764 3644 -19752
rect 4604 -19176 4662 -19164
rect 4604 -19752 4616 -19176
rect 4650 -19752 4662 -19176
rect 4604 -19764 4662 -19752
rect 5622 -19176 5680 -19164
rect 5622 -19752 5634 -19176
rect 5668 -19752 5680 -19176
rect 5622 -19764 5680 -19752
rect 6640 -19176 6698 -19164
rect 6640 -19752 6652 -19176
rect 6686 -19752 6698 -19176
rect 6640 -19764 6698 -19752
rect 7658 -19176 7716 -19164
rect 7658 -19752 7670 -19176
rect 7704 -19752 7716 -19176
rect 7658 -19764 7716 -19752
rect 8676 -19176 8734 -19164
rect 8676 -19752 8688 -19176
rect 8722 -19752 8734 -19176
rect 8676 -19764 8734 -19752
rect 9694 -19176 9752 -19164
rect 9694 -19752 9706 -19176
rect 9740 -19752 9752 -19176
rect 9694 -19764 9752 -19752
rect 10712 -19176 10770 -19164
rect 10712 -19752 10724 -19176
rect 10758 -19752 10770 -19176
rect 10712 -19764 10770 -19752
rect 11730 -19176 11788 -19164
rect 11730 -19752 11742 -19176
rect 11776 -19752 11788 -19176
rect 11730 -19764 11788 -19752
rect 12748 -19176 12806 -19164
rect 12748 -19752 12760 -19176
rect 12794 -19752 12806 -19176
rect 12748 -19764 12806 -19752
rect 13766 -19176 13824 -19164
rect 13766 -19752 13778 -19176
rect 13812 -19752 13824 -19176
rect 13766 -19764 13824 -19752
rect 14784 -19176 14842 -19164
rect 14784 -19752 14796 -19176
rect 14830 -19752 14842 -19176
rect 14784 -19764 14842 -19752
rect 15802 -19176 15860 -19164
rect 15802 -19752 15814 -19176
rect 15848 -19752 15860 -19176
rect 15802 -19764 15860 -19752
rect 16820 -19176 16878 -19164
rect 16820 -19752 16832 -19176
rect 16866 -19752 16878 -19176
rect 16820 -19764 16878 -19752
rect 17838 -19176 17896 -19164
rect 17838 -19752 17850 -19176
rect 17884 -19752 17896 -19176
rect 17838 -19764 17896 -19752
rect 18856 -19176 18914 -19164
rect 18856 -19752 18868 -19176
rect 18902 -19752 18914 -19176
rect 18856 -19764 18914 -19752
rect 19874 -19176 19932 -19164
rect 19874 -19752 19886 -19176
rect 19920 -19752 19932 -19176
rect 19874 -19764 19932 -19752
rect 20892 -19176 20950 -19164
rect 20892 -19752 20904 -19176
rect 20938 -19752 20950 -19176
rect 20892 -19764 20950 -19752
rect 21910 -19176 21968 -19164
rect 21910 -19752 21922 -19176
rect 21956 -19752 21968 -19176
rect 21910 -19764 21968 -19752
rect 22928 -19176 22986 -19164
rect 22928 -19752 22940 -19176
rect 22974 -19752 22986 -19176
rect 22928 -19764 22986 -19752
rect 2568 -20410 2626 -20398
rect 2568 -20986 2580 -20410
rect 2614 -20986 2626 -20410
rect 2568 -20998 2626 -20986
rect 3586 -20410 3644 -20398
rect 3586 -20986 3598 -20410
rect 3632 -20986 3644 -20410
rect 3586 -20998 3644 -20986
rect 4604 -20410 4662 -20398
rect 4604 -20986 4616 -20410
rect 4650 -20986 4662 -20410
rect 4604 -20998 4662 -20986
rect 5622 -20410 5680 -20398
rect 5622 -20986 5634 -20410
rect 5668 -20986 5680 -20410
rect 5622 -20998 5680 -20986
rect 6640 -20410 6698 -20398
rect 6640 -20986 6652 -20410
rect 6686 -20986 6698 -20410
rect 6640 -20998 6698 -20986
rect 7658 -20410 7716 -20398
rect 7658 -20986 7670 -20410
rect 7704 -20986 7716 -20410
rect 7658 -20998 7716 -20986
rect 8676 -20410 8734 -20398
rect 8676 -20986 8688 -20410
rect 8722 -20986 8734 -20410
rect 8676 -20998 8734 -20986
rect 9694 -20410 9752 -20398
rect 9694 -20986 9706 -20410
rect 9740 -20986 9752 -20410
rect 9694 -20998 9752 -20986
rect 10712 -20410 10770 -20398
rect 10712 -20986 10724 -20410
rect 10758 -20986 10770 -20410
rect 10712 -20998 10770 -20986
rect 11730 -20410 11788 -20398
rect 11730 -20986 11742 -20410
rect 11776 -20986 11788 -20410
rect 11730 -20998 11788 -20986
rect 12748 -20410 12806 -20398
rect 12748 -20986 12760 -20410
rect 12794 -20986 12806 -20410
rect 12748 -20998 12806 -20986
rect 13766 -20410 13824 -20398
rect 13766 -20986 13778 -20410
rect 13812 -20986 13824 -20410
rect 13766 -20998 13824 -20986
rect 14784 -20410 14842 -20398
rect 14784 -20986 14796 -20410
rect 14830 -20986 14842 -20410
rect 14784 -20998 14842 -20986
rect 15802 -20410 15860 -20398
rect 15802 -20986 15814 -20410
rect 15848 -20986 15860 -20410
rect 15802 -20998 15860 -20986
rect 16820 -20410 16878 -20398
rect 16820 -20986 16832 -20410
rect 16866 -20986 16878 -20410
rect 16820 -20998 16878 -20986
rect 17838 -20410 17896 -20398
rect 17838 -20986 17850 -20410
rect 17884 -20986 17896 -20410
rect 17838 -20998 17896 -20986
rect 18856 -20410 18914 -20398
rect 18856 -20986 18868 -20410
rect 18902 -20986 18914 -20410
rect 18856 -20998 18914 -20986
rect 19874 -20410 19932 -20398
rect 19874 -20986 19886 -20410
rect 19920 -20986 19932 -20410
rect 19874 -20998 19932 -20986
rect 20892 -20410 20950 -20398
rect 20892 -20986 20904 -20410
rect 20938 -20986 20950 -20410
rect 20892 -20998 20950 -20986
rect 21910 -20410 21968 -20398
rect 21910 -20986 21922 -20410
rect 21956 -20986 21968 -20410
rect 21910 -20998 21968 -20986
rect 22928 -20410 22986 -20398
rect 22928 -20986 22940 -20410
rect 22974 -20986 22986 -20410
rect 22928 -20998 22986 -20986
rect 2568 -21644 2626 -21632
rect 2568 -22220 2580 -21644
rect 2614 -22220 2626 -21644
rect 2568 -22232 2626 -22220
rect 3586 -21644 3644 -21632
rect 3586 -22220 3598 -21644
rect 3632 -22220 3644 -21644
rect 3586 -22232 3644 -22220
rect 4604 -21644 4662 -21632
rect 4604 -22220 4616 -21644
rect 4650 -22220 4662 -21644
rect 4604 -22232 4662 -22220
rect 5622 -21644 5680 -21632
rect 5622 -22220 5634 -21644
rect 5668 -22220 5680 -21644
rect 5622 -22232 5680 -22220
rect 6640 -21644 6698 -21632
rect 6640 -22220 6652 -21644
rect 6686 -22220 6698 -21644
rect 6640 -22232 6698 -22220
rect 7658 -21644 7716 -21632
rect 7658 -22220 7670 -21644
rect 7704 -22220 7716 -21644
rect 7658 -22232 7716 -22220
rect 8676 -21644 8734 -21632
rect 8676 -22220 8688 -21644
rect 8722 -22220 8734 -21644
rect 8676 -22232 8734 -22220
rect 9694 -21644 9752 -21632
rect 9694 -22220 9706 -21644
rect 9740 -22220 9752 -21644
rect 9694 -22232 9752 -22220
rect 10712 -21644 10770 -21632
rect 10712 -22220 10724 -21644
rect 10758 -22220 10770 -21644
rect 10712 -22232 10770 -22220
rect 11730 -21644 11788 -21632
rect 11730 -22220 11742 -21644
rect 11776 -22220 11788 -21644
rect 11730 -22232 11788 -22220
rect 12748 -21644 12806 -21632
rect 12748 -22220 12760 -21644
rect 12794 -22220 12806 -21644
rect 12748 -22232 12806 -22220
rect 13766 -21644 13824 -21632
rect 13766 -22220 13778 -21644
rect 13812 -22220 13824 -21644
rect 13766 -22232 13824 -22220
rect 14784 -21644 14842 -21632
rect 14784 -22220 14796 -21644
rect 14830 -22220 14842 -21644
rect 14784 -22232 14842 -22220
rect 15802 -21644 15860 -21632
rect 15802 -22220 15814 -21644
rect 15848 -22220 15860 -21644
rect 15802 -22232 15860 -22220
rect 16820 -21644 16878 -21632
rect 16820 -22220 16832 -21644
rect 16866 -22220 16878 -21644
rect 16820 -22232 16878 -22220
rect 17838 -21644 17896 -21632
rect 17838 -22220 17850 -21644
rect 17884 -22220 17896 -21644
rect 17838 -22232 17896 -22220
rect 18856 -21644 18914 -21632
rect 18856 -22220 18868 -21644
rect 18902 -22220 18914 -21644
rect 18856 -22232 18914 -22220
rect 19874 -21644 19932 -21632
rect 19874 -22220 19886 -21644
rect 19920 -22220 19932 -21644
rect 19874 -22232 19932 -22220
rect 20892 -21644 20950 -21632
rect 20892 -22220 20904 -21644
rect 20938 -22220 20950 -21644
rect 20892 -22232 20950 -22220
rect 21910 -21644 21968 -21632
rect 21910 -22220 21922 -21644
rect 21956 -22220 21968 -21644
rect 21910 -22232 21968 -22220
rect 22928 -21644 22986 -21632
rect 22928 -22220 22940 -21644
rect 22974 -22220 22986 -21644
rect 22928 -22232 22986 -22220
rect 2568 -22876 2626 -22864
rect 2568 -23452 2580 -22876
rect 2614 -23452 2626 -22876
rect 2568 -23464 2626 -23452
rect 3586 -22876 3644 -22864
rect 3586 -23452 3598 -22876
rect 3632 -23452 3644 -22876
rect 3586 -23464 3644 -23452
rect 4604 -22876 4662 -22864
rect 4604 -23452 4616 -22876
rect 4650 -23452 4662 -22876
rect 4604 -23464 4662 -23452
rect 5622 -22876 5680 -22864
rect 5622 -23452 5634 -22876
rect 5668 -23452 5680 -22876
rect 5622 -23464 5680 -23452
rect 6640 -22876 6698 -22864
rect 6640 -23452 6652 -22876
rect 6686 -23452 6698 -22876
rect 6640 -23464 6698 -23452
rect 7658 -22876 7716 -22864
rect 7658 -23452 7670 -22876
rect 7704 -23452 7716 -22876
rect 7658 -23464 7716 -23452
rect 8676 -22876 8734 -22864
rect 8676 -23452 8688 -22876
rect 8722 -23452 8734 -22876
rect 8676 -23464 8734 -23452
rect 9694 -22876 9752 -22864
rect 9694 -23452 9706 -22876
rect 9740 -23452 9752 -22876
rect 9694 -23464 9752 -23452
rect 10712 -22876 10770 -22864
rect 10712 -23452 10724 -22876
rect 10758 -23452 10770 -22876
rect 10712 -23464 10770 -23452
rect 11730 -22876 11788 -22864
rect 11730 -23452 11742 -22876
rect 11776 -23452 11788 -22876
rect 11730 -23464 11788 -23452
rect 12748 -22876 12806 -22864
rect 12748 -23452 12760 -22876
rect 12794 -23452 12806 -22876
rect 12748 -23464 12806 -23452
rect 13766 -22876 13824 -22864
rect 13766 -23452 13778 -22876
rect 13812 -23452 13824 -22876
rect 13766 -23464 13824 -23452
rect 14784 -22876 14842 -22864
rect 14784 -23452 14796 -22876
rect 14830 -23452 14842 -22876
rect 14784 -23464 14842 -23452
rect 15802 -22876 15860 -22864
rect 15802 -23452 15814 -22876
rect 15848 -23452 15860 -22876
rect 15802 -23464 15860 -23452
rect 16820 -22876 16878 -22864
rect 16820 -23452 16832 -22876
rect 16866 -23452 16878 -22876
rect 16820 -23464 16878 -23452
rect 17838 -22876 17896 -22864
rect 17838 -23452 17850 -22876
rect 17884 -23452 17896 -22876
rect 17838 -23464 17896 -23452
rect 18856 -22876 18914 -22864
rect 18856 -23452 18868 -22876
rect 18902 -23452 18914 -22876
rect 18856 -23464 18914 -23452
rect 19874 -22876 19932 -22864
rect 19874 -23452 19886 -22876
rect 19920 -23452 19932 -22876
rect 19874 -23464 19932 -23452
rect 20892 -22876 20950 -22864
rect 20892 -23452 20904 -22876
rect 20938 -23452 20950 -22876
rect 20892 -23464 20950 -23452
rect 21910 -22876 21968 -22864
rect 21910 -23452 21922 -22876
rect 21956 -23452 21968 -22876
rect 21910 -23464 21968 -23452
rect 22928 -22876 22986 -22864
rect 22928 -23452 22940 -22876
rect 22974 -23452 22986 -22876
rect 22928 -23464 22986 -23452
rect 2568 -24110 2626 -24098
rect 2568 -24686 2580 -24110
rect 2614 -24686 2626 -24110
rect 2568 -24698 2626 -24686
rect 3586 -24110 3644 -24098
rect 3586 -24686 3598 -24110
rect 3632 -24686 3644 -24110
rect 3586 -24698 3644 -24686
rect 4604 -24110 4662 -24098
rect 4604 -24686 4616 -24110
rect 4650 -24686 4662 -24110
rect 4604 -24698 4662 -24686
rect 5622 -24110 5680 -24098
rect 5622 -24686 5634 -24110
rect 5668 -24686 5680 -24110
rect 5622 -24698 5680 -24686
rect 6640 -24110 6698 -24098
rect 6640 -24686 6652 -24110
rect 6686 -24686 6698 -24110
rect 6640 -24698 6698 -24686
rect 7658 -24110 7716 -24098
rect 7658 -24686 7670 -24110
rect 7704 -24686 7716 -24110
rect 7658 -24698 7716 -24686
rect 8676 -24110 8734 -24098
rect 8676 -24686 8688 -24110
rect 8722 -24686 8734 -24110
rect 8676 -24698 8734 -24686
rect 9694 -24110 9752 -24098
rect 9694 -24686 9706 -24110
rect 9740 -24686 9752 -24110
rect 9694 -24698 9752 -24686
rect 10712 -24110 10770 -24098
rect 10712 -24686 10724 -24110
rect 10758 -24686 10770 -24110
rect 10712 -24698 10770 -24686
rect 11730 -24110 11788 -24098
rect 11730 -24686 11742 -24110
rect 11776 -24686 11788 -24110
rect 11730 -24698 11788 -24686
rect 12748 -24110 12806 -24098
rect 12748 -24686 12760 -24110
rect 12794 -24686 12806 -24110
rect 12748 -24698 12806 -24686
rect 13766 -24110 13824 -24098
rect 13766 -24686 13778 -24110
rect 13812 -24686 13824 -24110
rect 13766 -24698 13824 -24686
rect 14784 -24110 14842 -24098
rect 14784 -24686 14796 -24110
rect 14830 -24686 14842 -24110
rect 14784 -24698 14842 -24686
rect 15802 -24110 15860 -24098
rect 15802 -24686 15814 -24110
rect 15848 -24686 15860 -24110
rect 15802 -24698 15860 -24686
rect 16820 -24110 16878 -24098
rect 16820 -24686 16832 -24110
rect 16866 -24686 16878 -24110
rect 16820 -24698 16878 -24686
rect 17838 -24110 17896 -24098
rect 17838 -24686 17850 -24110
rect 17884 -24686 17896 -24110
rect 17838 -24698 17896 -24686
rect 18856 -24110 18914 -24098
rect 18856 -24686 18868 -24110
rect 18902 -24686 18914 -24110
rect 18856 -24698 18914 -24686
rect 19874 -24110 19932 -24098
rect 19874 -24686 19886 -24110
rect 19920 -24686 19932 -24110
rect 19874 -24698 19932 -24686
rect 20892 -24110 20950 -24098
rect 20892 -24686 20904 -24110
rect 20938 -24686 20950 -24110
rect 20892 -24698 20950 -24686
rect 21910 -24110 21968 -24098
rect 21910 -24686 21922 -24110
rect 21956 -24686 21968 -24110
rect 21910 -24698 21968 -24686
rect 22928 -24110 22986 -24098
rect 22928 -24686 22940 -24110
rect 22974 -24686 22986 -24110
rect 22928 -24698 22986 -24686
<< ndiffc >>
rect -9184 -13100 -9150 -12524
rect -8166 -13100 -8132 -12524
rect -7148 -13100 -7114 -12524
rect -6130 -13100 -6096 -12524
rect -5112 -13100 -5078 -12524
rect -4094 -13100 -4060 -12524
rect -3076 -13100 -3042 -12524
rect -2058 -13100 -2024 -12524
rect -1040 -13100 -1006 -12524
rect -22 -13100 12 -12524
rect -9184 -13918 -9150 -13342
rect -8166 -13918 -8132 -13342
rect -7148 -13918 -7114 -13342
rect -6130 -13918 -6096 -13342
rect -5112 -13918 -5078 -13342
rect -4094 -13918 -4060 -13342
rect -3076 -13918 -3042 -13342
rect -2058 -13918 -2024 -13342
rect -1040 -13918 -1006 -13342
rect -22 -13918 12 -13342
rect -9184 -14736 -9150 -14160
rect -8166 -14736 -8132 -14160
rect -7148 -14736 -7114 -14160
rect -6130 -14736 -6096 -14160
rect -5112 -14736 -5078 -14160
rect -4094 -14736 -4060 -14160
rect -3076 -14736 -3042 -14160
rect -2058 -14736 -2024 -14160
rect -1040 -14736 -1006 -14160
rect -22 -14736 12 -14160
rect 2582 -14820 2616 -14244
rect 3600 -14820 3634 -14244
rect 4618 -14820 4652 -14244
rect 5636 -14820 5670 -14244
rect 6654 -14820 6688 -14244
rect 7672 -14820 7706 -14244
rect 8690 -14820 8724 -14244
rect 9708 -14820 9742 -14244
rect 10726 -14820 10760 -14244
rect 11744 -14820 11778 -14244
rect 12762 -14820 12796 -14244
rect 13780 -14820 13814 -14244
rect 14798 -14820 14832 -14244
rect 15816 -14820 15850 -14244
rect 16834 -14820 16868 -14244
rect 17852 -14820 17886 -14244
rect 18870 -14820 18904 -14244
rect 19888 -14820 19922 -14244
rect 20906 -14820 20940 -14244
rect 21924 -14820 21958 -14244
rect 22942 -14820 22976 -14244
rect -9184 -15554 -9150 -14978
rect -8166 -15554 -8132 -14978
rect -7148 -15554 -7114 -14978
rect -6130 -15554 -6096 -14978
rect -5112 -15554 -5078 -14978
rect -4094 -15554 -4060 -14978
rect -3076 -15554 -3042 -14978
rect -2058 -15554 -2024 -14978
rect -1040 -15554 -1006 -14978
rect -22 -15554 12 -14978
rect -9184 -16372 -9150 -15796
rect -8166 -16372 -8132 -15796
rect -7148 -16372 -7114 -15796
rect -6130 -16372 -6096 -15796
rect -5112 -16372 -5078 -15796
rect -4094 -16372 -4060 -15796
rect -3076 -16372 -3042 -15796
rect -2058 -16372 -2024 -15796
rect -1040 -16372 -1006 -15796
rect -22 -16372 12 -15796
rect 2582 -16052 2616 -15476
rect 3600 -16052 3634 -15476
rect 4618 -16052 4652 -15476
rect 5636 -16052 5670 -15476
rect 6654 -16052 6688 -15476
rect 7672 -16052 7706 -15476
rect 8690 -16052 8724 -15476
rect 9708 -16052 9742 -15476
rect 10726 -16052 10760 -15476
rect 11744 -16052 11778 -15476
rect 12762 -16052 12796 -15476
rect 13780 -16052 13814 -15476
rect 14798 -16052 14832 -15476
rect 15816 -16052 15850 -15476
rect 16834 -16052 16868 -15476
rect 17852 -16052 17886 -15476
rect 18870 -16052 18904 -15476
rect 19888 -16052 19922 -15476
rect 20906 -16052 20940 -15476
rect 21924 -16052 21958 -15476
rect 22942 -16052 22976 -15476
rect -9184 -17190 -9150 -16614
rect -8166 -17190 -8132 -16614
rect -7148 -17190 -7114 -16614
rect -6130 -17190 -6096 -16614
rect -5112 -17190 -5078 -16614
rect -4094 -17190 -4060 -16614
rect -3076 -17190 -3042 -16614
rect -2058 -17190 -2024 -16614
rect -1040 -17190 -1006 -16614
rect -22 -17190 12 -16614
rect 2580 -17286 2614 -16710
rect 3598 -17286 3632 -16710
rect 4616 -17286 4650 -16710
rect 5634 -17286 5668 -16710
rect 6652 -17286 6686 -16710
rect 7670 -17286 7704 -16710
rect 8688 -17286 8722 -16710
rect 9706 -17286 9740 -16710
rect 10724 -17286 10758 -16710
rect 11742 -17286 11776 -16710
rect 12760 -17286 12794 -16710
rect 13778 -17286 13812 -16710
rect 14796 -17286 14830 -16710
rect 15814 -17286 15848 -16710
rect 16832 -17286 16866 -16710
rect 17850 -17286 17884 -16710
rect 18868 -17286 18902 -16710
rect 19886 -17286 19920 -16710
rect 20904 -17286 20938 -16710
rect 21922 -17286 21956 -16710
rect 22940 -17286 22974 -16710
rect -9184 -18008 -9150 -17432
rect -8166 -18008 -8132 -17432
rect -7148 -18008 -7114 -17432
rect -6130 -18008 -6096 -17432
rect -5112 -18008 -5078 -17432
rect -4094 -18008 -4060 -17432
rect -3076 -18008 -3042 -17432
rect -2058 -18008 -2024 -17432
rect -1040 -18008 -1006 -17432
rect -22 -18008 12 -17432
rect -9184 -18826 -9150 -18250
rect -8166 -18826 -8132 -18250
rect -7148 -18826 -7114 -18250
rect -6130 -18826 -6096 -18250
rect -5112 -18826 -5078 -18250
rect -4094 -18826 -4060 -18250
rect -3076 -18826 -3042 -18250
rect -2058 -18826 -2024 -18250
rect -1040 -18826 -1006 -18250
rect -22 -18826 12 -18250
rect 2580 -18520 2614 -17944
rect 3598 -18520 3632 -17944
rect 4616 -18520 4650 -17944
rect 5634 -18520 5668 -17944
rect 6652 -18520 6686 -17944
rect 7670 -18520 7704 -17944
rect 8688 -18520 8722 -17944
rect 9706 -18520 9740 -17944
rect 10724 -18520 10758 -17944
rect 11742 -18520 11776 -17944
rect 12760 -18520 12794 -17944
rect 13778 -18520 13812 -17944
rect 14796 -18520 14830 -17944
rect 15814 -18520 15848 -17944
rect 16832 -18520 16866 -17944
rect 17850 -18520 17884 -17944
rect 18868 -18520 18902 -17944
rect 19886 -18520 19920 -17944
rect 20904 -18520 20938 -17944
rect 21922 -18520 21956 -17944
rect 22940 -18520 22974 -17944
rect 2580 -19752 2614 -19176
rect 3598 -19752 3632 -19176
rect 4616 -19752 4650 -19176
rect 5634 -19752 5668 -19176
rect 6652 -19752 6686 -19176
rect 7670 -19752 7704 -19176
rect 8688 -19752 8722 -19176
rect 9706 -19752 9740 -19176
rect 10724 -19752 10758 -19176
rect 11742 -19752 11776 -19176
rect 12760 -19752 12794 -19176
rect 13778 -19752 13812 -19176
rect 14796 -19752 14830 -19176
rect 15814 -19752 15848 -19176
rect 16832 -19752 16866 -19176
rect 17850 -19752 17884 -19176
rect 18868 -19752 18902 -19176
rect 19886 -19752 19920 -19176
rect 20904 -19752 20938 -19176
rect 21922 -19752 21956 -19176
rect 22940 -19752 22974 -19176
rect 2580 -20986 2614 -20410
rect 3598 -20986 3632 -20410
rect 4616 -20986 4650 -20410
rect 5634 -20986 5668 -20410
rect 6652 -20986 6686 -20410
rect 7670 -20986 7704 -20410
rect 8688 -20986 8722 -20410
rect 9706 -20986 9740 -20410
rect 10724 -20986 10758 -20410
rect 11742 -20986 11776 -20410
rect 12760 -20986 12794 -20410
rect 13778 -20986 13812 -20410
rect 14796 -20986 14830 -20410
rect 15814 -20986 15848 -20410
rect 16832 -20986 16866 -20410
rect 17850 -20986 17884 -20410
rect 18868 -20986 18902 -20410
rect 19886 -20986 19920 -20410
rect 20904 -20986 20938 -20410
rect 21922 -20986 21956 -20410
rect 22940 -20986 22974 -20410
rect 2580 -22220 2614 -21644
rect 3598 -22220 3632 -21644
rect 4616 -22220 4650 -21644
rect 5634 -22220 5668 -21644
rect 6652 -22220 6686 -21644
rect 7670 -22220 7704 -21644
rect 8688 -22220 8722 -21644
rect 9706 -22220 9740 -21644
rect 10724 -22220 10758 -21644
rect 11742 -22220 11776 -21644
rect 12760 -22220 12794 -21644
rect 13778 -22220 13812 -21644
rect 14796 -22220 14830 -21644
rect 15814 -22220 15848 -21644
rect 16832 -22220 16866 -21644
rect 17850 -22220 17884 -21644
rect 18868 -22220 18902 -21644
rect 19886 -22220 19920 -21644
rect 20904 -22220 20938 -21644
rect 21922 -22220 21956 -21644
rect 22940 -22220 22974 -21644
rect 2580 -23452 2614 -22876
rect 3598 -23452 3632 -22876
rect 4616 -23452 4650 -22876
rect 5634 -23452 5668 -22876
rect 6652 -23452 6686 -22876
rect 7670 -23452 7704 -22876
rect 8688 -23452 8722 -22876
rect 9706 -23452 9740 -22876
rect 10724 -23452 10758 -22876
rect 11742 -23452 11776 -22876
rect 12760 -23452 12794 -22876
rect 13778 -23452 13812 -22876
rect 14796 -23452 14830 -22876
rect 15814 -23452 15848 -22876
rect 16832 -23452 16866 -22876
rect 17850 -23452 17884 -22876
rect 18868 -23452 18902 -22876
rect 19886 -23452 19920 -22876
rect 20904 -23452 20938 -22876
rect 21922 -23452 21956 -22876
rect 22940 -23452 22974 -22876
rect 2580 -24686 2614 -24110
rect 3598 -24686 3632 -24110
rect 4616 -24686 4650 -24110
rect 5634 -24686 5668 -24110
rect 6652 -24686 6686 -24110
rect 7670 -24686 7704 -24110
rect 8688 -24686 8722 -24110
rect 9706 -24686 9740 -24110
rect 10724 -24686 10758 -24110
rect 11742 -24686 11776 -24110
rect 12760 -24686 12794 -24110
rect 13778 -24686 13812 -24110
rect 14796 -24686 14830 -24110
rect 15814 -24686 15848 -24110
rect 16832 -24686 16866 -24110
rect 17850 -24686 17884 -24110
rect 18868 -24686 18902 -24110
rect 19886 -24686 19920 -24110
rect 20904 -24686 20938 -24110
rect 21922 -24686 21956 -24110
rect 22940 -24686 22974 -24110
<< psubdiff >>
rect -12322 -11278 -12160 -11178
rect 24760 -11278 24922 -11178
rect -12322 -11340 -12222 -11278
rect 24822 -11340 24922 -11278
rect -12322 -27122 -12222 -27060
rect 24822 -27122 24922 -27060
rect -12322 -27222 -12160 -27122
rect 24760 -27222 24922 -27122
<< nsubdiff >>
rect 378 4222 540 4322
rect 24660 4222 24822 4322
rect 378 4160 478 4222
rect 378 -10248 478 -10186
rect 24722 4160 24822 4222
rect 24722 -10248 24822 -10186
rect 378 -10348 540 -10248
rect 24660 -10348 24822 -10248
<< psubdiffcont >>
rect -12160 -11278 24760 -11178
rect -12322 -27060 -12222 -11340
rect 24822 -27060 24922 -11340
rect -12160 -27222 24760 -27122
<< nsubdiffcont >>
rect 540 4222 24660 4322
rect 378 -10186 478 4160
rect 24722 -10186 24822 4160
rect 540 -10348 24660 -10248
<< poly >>
rect -8952 -12440 -8364 -12424
rect -8952 -12457 -8936 -12440
rect -9138 -12474 -8936 -12457
rect -8380 -12457 -8364 -12440
rect -7934 -12440 -7346 -12424
rect -7934 -12457 -7918 -12440
rect -8380 -12474 -8178 -12457
rect -9138 -12512 -8178 -12474
rect -8120 -12474 -7918 -12457
rect -7362 -12457 -7346 -12440
rect -6916 -12440 -6328 -12424
rect -6916 -12457 -6900 -12440
rect -7362 -12474 -7160 -12457
rect -8120 -12512 -7160 -12474
rect -7102 -12474 -6900 -12457
rect -6344 -12457 -6328 -12440
rect -5898 -12440 -5310 -12424
rect -5898 -12457 -5882 -12440
rect -6344 -12474 -6142 -12457
rect -7102 -12512 -6142 -12474
rect -6084 -12474 -5882 -12457
rect -5326 -12457 -5310 -12440
rect -4880 -12440 -4292 -12424
rect -4880 -12457 -4864 -12440
rect -5326 -12474 -5124 -12457
rect -6084 -12512 -5124 -12474
rect -5066 -12474 -4864 -12457
rect -4308 -12457 -4292 -12440
rect -3862 -12440 -3274 -12424
rect -3862 -12457 -3846 -12440
rect -4308 -12474 -4106 -12457
rect -5066 -12512 -4106 -12474
rect -4048 -12474 -3846 -12457
rect -3290 -12457 -3274 -12440
rect -2844 -12440 -2256 -12424
rect -2844 -12457 -2828 -12440
rect -3290 -12474 -3088 -12457
rect -4048 -12512 -3088 -12474
rect -3030 -12474 -2828 -12457
rect -2272 -12457 -2256 -12440
rect -1826 -12440 -1238 -12424
rect -1826 -12457 -1810 -12440
rect -2272 -12474 -2070 -12457
rect -3030 -12512 -2070 -12474
rect -2012 -12474 -1810 -12457
rect -1254 -12457 -1238 -12440
rect -808 -12440 -220 -12424
rect -808 -12457 -792 -12440
rect -1254 -12474 -1052 -12457
rect -2012 -12512 -1052 -12474
rect -994 -12474 -792 -12457
rect -236 -12457 -220 -12440
rect -236 -12474 -34 -12457
rect -994 -12512 -34 -12474
rect -9138 -13150 -8178 -13112
rect -9138 -13167 -8936 -13150
rect -8952 -13184 -8936 -13167
rect -8380 -13167 -8178 -13150
rect -8120 -13150 -7160 -13112
rect -8120 -13167 -7918 -13150
rect -8380 -13184 -8364 -13167
rect -8952 -13200 -8364 -13184
rect -7934 -13184 -7918 -13167
rect -7362 -13167 -7160 -13150
rect -7102 -13150 -6142 -13112
rect -7102 -13167 -6900 -13150
rect -7362 -13184 -7346 -13167
rect -7934 -13200 -7346 -13184
rect -6916 -13184 -6900 -13167
rect -6344 -13167 -6142 -13150
rect -6084 -13150 -5124 -13112
rect -6084 -13167 -5882 -13150
rect -6344 -13184 -6328 -13167
rect -6916 -13200 -6328 -13184
rect -5898 -13184 -5882 -13167
rect -5326 -13167 -5124 -13150
rect -5066 -13150 -4106 -13112
rect -5066 -13167 -4864 -13150
rect -5326 -13184 -5310 -13167
rect -5898 -13200 -5310 -13184
rect -4880 -13184 -4864 -13167
rect -4308 -13167 -4106 -13150
rect -4048 -13150 -3088 -13112
rect -4048 -13167 -3846 -13150
rect -4308 -13184 -4292 -13167
rect -4880 -13200 -4292 -13184
rect -3862 -13184 -3846 -13167
rect -3290 -13167 -3088 -13150
rect -3030 -13150 -2070 -13112
rect -3030 -13167 -2828 -13150
rect -3290 -13184 -3274 -13167
rect -3862 -13200 -3274 -13184
rect -2844 -13184 -2828 -13167
rect -2272 -13167 -2070 -13150
rect -2012 -13150 -1052 -13112
rect -2012 -13167 -1810 -13150
rect -2272 -13184 -2256 -13167
rect -2844 -13200 -2256 -13184
rect -1826 -13184 -1810 -13167
rect -1254 -13167 -1052 -13150
rect -994 -13150 -34 -13112
rect -994 -13167 -792 -13150
rect -1254 -13184 -1238 -13167
rect -1826 -13200 -1238 -13184
rect -808 -13184 -792 -13167
rect -236 -13167 -34 -13150
rect -236 -13184 -220 -13167
rect -808 -13200 -220 -13184
rect -8952 -13258 -8364 -13242
rect -8952 -13275 -8936 -13258
rect -9138 -13292 -8936 -13275
rect -8380 -13275 -8364 -13258
rect -7934 -13258 -7346 -13242
rect -7934 -13275 -7918 -13258
rect -8380 -13292 -8178 -13275
rect -9138 -13330 -8178 -13292
rect -8120 -13292 -7918 -13275
rect -7362 -13275 -7346 -13258
rect -6916 -13258 -6328 -13242
rect -6916 -13275 -6900 -13258
rect -7362 -13292 -7160 -13275
rect -8120 -13330 -7160 -13292
rect -7102 -13292 -6900 -13275
rect -6344 -13275 -6328 -13258
rect -5898 -13258 -5310 -13242
rect -5898 -13275 -5882 -13258
rect -6344 -13292 -6142 -13275
rect -7102 -13330 -6142 -13292
rect -6084 -13292 -5882 -13275
rect -5326 -13275 -5310 -13258
rect -4880 -13258 -4292 -13242
rect -4880 -13275 -4864 -13258
rect -5326 -13292 -5124 -13275
rect -6084 -13330 -5124 -13292
rect -5066 -13292 -4864 -13275
rect -4308 -13275 -4292 -13258
rect -3862 -13258 -3274 -13242
rect -3862 -13275 -3846 -13258
rect -4308 -13292 -4106 -13275
rect -5066 -13330 -4106 -13292
rect -4048 -13292 -3846 -13275
rect -3290 -13275 -3274 -13258
rect -2844 -13258 -2256 -13242
rect -2844 -13275 -2828 -13258
rect -3290 -13292 -3088 -13275
rect -4048 -13330 -3088 -13292
rect -3030 -13292 -2828 -13275
rect -2272 -13275 -2256 -13258
rect -1826 -13258 -1238 -13242
rect -1826 -13275 -1810 -13258
rect -2272 -13292 -2070 -13275
rect -3030 -13330 -2070 -13292
rect -2012 -13292 -1810 -13275
rect -1254 -13275 -1238 -13258
rect -808 -13258 -220 -13242
rect -808 -13275 -792 -13258
rect -1254 -13292 -1052 -13275
rect -2012 -13330 -1052 -13292
rect -994 -13292 -792 -13275
rect -236 -13275 -220 -13258
rect -236 -13292 -34 -13275
rect -994 -13330 -34 -13292
rect -9138 -13968 -8178 -13930
rect -9138 -13985 -8936 -13968
rect -8952 -14002 -8936 -13985
rect -8380 -13985 -8178 -13968
rect -8120 -13968 -7160 -13930
rect -8120 -13985 -7918 -13968
rect -8380 -14002 -8364 -13985
rect -8952 -14018 -8364 -14002
rect -7934 -14002 -7918 -13985
rect -7362 -13985 -7160 -13968
rect -7102 -13968 -6142 -13930
rect -7102 -13985 -6900 -13968
rect -7362 -14002 -7346 -13985
rect -7934 -14018 -7346 -14002
rect -6916 -14002 -6900 -13985
rect -6344 -13985 -6142 -13968
rect -6084 -13968 -5124 -13930
rect -6084 -13985 -5882 -13968
rect -6344 -14002 -6328 -13985
rect -6916 -14018 -6328 -14002
rect -5898 -14002 -5882 -13985
rect -5326 -13985 -5124 -13968
rect -5066 -13968 -4106 -13930
rect -5066 -13985 -4864 -13968
rect -5326 -14002 -5310 -13985
rect -5898 -14018 -5310 -14002
rect -4880 -14002 -4864 -13985
rect -4308 -13985 -4106 -13968
rect -4048 -13968 -3088 -13930
rect -4048 -13985 -3846 -13968
rect -4308 -14002 -4292 -13985
rect -4880 -14018 -4292 -14002
rect -3862 -14002 -3846 -13985
rect -3290 -13985 -3088 -13968
rect -3030 -13968 -2070 -13930
rect -3030 -13985 -2828 -13968
rect -3290 -14002 -3274 -13985
rect -3862 -14018 -3274 -14002
rect -2844 -14002 -2828 -13985
rect -2272 -13985 -2070 -13968
rect -2012 -13968 -1052 -13930
rect -2012 -13985 -1810 -13968
rect -2272 -14002 -2256 -13985
rect -2844 -14018 -2256 -14002
rect -1826 -14002 -1810 -13985
rect -1254 -13985 -1052 -13968
rect -994 -13968 -34 -13930
rect -994 -13985 -792 -13968
rect -1254 -14002 -1238 -13985
rect -1826 -14018 -1238 -14002
rect -808 -14002 -792 -13985
rect -236 -13985 -34 -13968
rect -236 -14002 -220 -13985
rect -808 -14018 -220 -14002
rect -8952 -14076 -8364 -14060
rect -8952 -14093 -8936 -14076
rect -9138 -14110 -8936 -14093
rect -8380 -14093 -8364 -14076
rect -7934 -14076 -7346 -14060
rect -7934 -14093 -7918 -14076
rect -8380 -14110 -8178 -14093
rect -9138 -14148 -8178 -14110
rect -8120 -14110 -7918 -14093
rect -7362 -14093 -7346 -14076
rect -6916 -14076 -6328 -14060
rect -6916 -14093 -6900 -14076
rect -7362 -14110 -7160 -14093
rect -8120 -14148 -7160 -14110
rect -7102 -14110 -6900 -14093
rect -6344 -14093 -6328 -14076
rect -5898 -14076 -5310 -14060
rect -5898 -14093 -5882 -14076
rect -6344 -14110 -6142 -14093
rect -7102 -14148 -6142 -14110
rect -6084 -14110 -5882 -14093
rect -5326 -14093 -5310 -14076
rect -4880 -14076 -4292 -14060
rect -4880 -14093 -4864 -14076
rect -5326 -14110 -5124 -14093
rect -6084 -14148 -5124 -14110
rect -5066 -14110 -4864 -14093
rect -4308 -14093 -4292 -14076
rect -3862 -14076 -3274 -14060
rect -3862 -14093 -3846 -14076
rect -4308 -14110 -4106 -14093
rect -5066 -14148 -4106 -14110
rect -4048 -14110 -3846 -14093
rect -3290 -14093 -3274 -14076
rect -2844 -14076 -2256 -14060
rect -2844 -14093 -2828 -14076
rect -3290 -14110 -3088 -14093
rect -4048 -14148 -3088 -14110
rect -3030 -14110 -2828 -14093
rect -2272 -14093 -2256 -14076
rect -1826 -14076 -1238 -14060
rect -1826 -14093 -1810 -14076
rect -2272 -14110 -2070 -14093
rect -3030 -14148 -2070 -14110
rect -2012 -14110 -1810 -14093
rect -1254 -14093 -1238 -14076
rect -808 -14076 -220 -14060
rect -808 -14093 -792 -14076
rect -1254 -14110 -1052 -14093
rect -2012 -14148 -1052 -14110
rect -994 -14110 -792 -14093
rect -236 -14093 -220 -14076
rect -236 -14110 -34 -14093
rect -994 -14148 -34 -14110
rect 2814 -14160 3402 -14144
rect 2814 -14177 2830 -14160
rect 2628 -14194 2830 -14177
rect 3386 -14177 3402 -14160
rect 3832 -14160 4420 -14144
rect 3832 -14177 3848 -14160
rect 3386 -14194 3588 -14177
rect 2628 -14232 3588 -14194
rect 3646 -14194 3848 -14177
rect 4404 -14177 4420 -14160
rect 4850 -14160 5438 -14144
rect 4850 -14177 4866 -14160
rect 4404 -14194 4606 -14177
rect 3646 -14232 4606 -14194
rect 4664 -14194 4866 -14177
rect 5422 -14177 5438 -14160
rect 5868 -14160 6456 -14144
rect 5868 -14177 5884 -14160
rect 5422 -14194 5624 -14177
rect 4664 -14232 5624 -14194
rect 5682 -14194 5884 -14177
rect 6440 -14177 6456 -14160
rect 6886 -14160 7474 -14144
rect 6886 -14177 6902 -14160
rect 6440 -14194 6642 -14177
rect 5682 -14232 6642 -14194
rect 6700 -14194 6902 -14177
rect 7458 -14177 7474 -14160
rect 7904 -14160 8492 -14144
rect 7904 -14177 7920 -14160
rect 7458 -14194 7660 -14177
rect 6700 -14232 7660 -14194
rect 7718 -14194 7920 -14177
rect 8476 -14177 8492 -14160
rect 8922 -14160 9510 -14144
rect 8922 -14177 8938 -14160
rect 8476 -14194 8678 -14177
rect 7718 -14232 8678 -14194
rect 8736 -14194 8938 -14177
rect 9494 -14177 9510 -14160
rect 9940 -14160 10528 -14144
rect 9940 -14177 9956 -14160
rect 9494 -14194 9696 -14177
rect 8736 -14232 9696 -14194
rect 9754 -14194 9956 -14177
rect 10512 -14177 10528 -14160
rect 10958 -14160 11546 -14144
rect 10958 -14177 10974 -14160
rect 10512 -14194 10714 -14177
rect 9754 -14232 10714 -14194
rect 10772 -14194 10974 -14177
rect 11530 -14177 11546 -14160
rect 11976 -14160 12564 -14144
rect 11976 -14177 11992 -14160
rect 11530 -14194 11732 -14177
rect 10772 -14232 11732 -14194
rect 11790 -14194 11992 -14177
rect 12548 -14177 12564 -14160
rect 12994 -14160 13582 -14144
rect 12994 -14177 13010 -14160
rect 12548 -14194 12750 -14177
rect 11790 -14232 12750 -14194
rect 12808 -14194 13010 -14177
rect 13566 -14177 13582 -14160
rect 14012 -14160 14600 -14144
rect 14012 -14177 14028 -14160
rect 13566 -14194 13768 -14177
rect 12808 -14232 13768 -14194
rect 13826 -14194 14028 -14177
rect 14584 -14177 14600 -14160
rect 15030 -14160 15618 -14144
rect 15030 -14177 15046 -14160
rect 14584 -14194 14786 -14177
rect 13826 -14232 14786 -14194
rect 14844 -14194 15046 -14177
rect 15602 -14177 15618 -14160
rect 16048 -14160 16636 -14144
rect 16048 -14177 16064 -14160
rect 15602 -14194 15804 -14177
rect 14844 -14232 15804 -14194
rect 15862 -14194 16064 -14177
rect 16620 -14177 16636 -14160
rect 17066 -14160 17654 -14144
rect 17066 -14177 17082 -14160
rect 16620 -14194 16822 -14177
rect 15862 -14232 16822 -14194
rect 16880 -14194 17082 -14177
rect 17638 -14177 17654 -14160
rect 18084 -14160 18672 -14144
rect 18084 -14177 18100 -14160
rect 17638 -14194 17840 -14177
rect 16880 -14232 17840 -14194
rect 17898 -14194 18100 -14177
rect 18656 -14177 18672 -14160
rect 19102 -14160 19690 -14144
rect 19102 -14177 19118 -14160
rect 18656 -14194 18858 -14177
rect 17898 -14232 18858 -14194
rect 18916 -14194 19118 -14177
rect 19674 -14177 19690 -14160
rect 20120 -14160 20708 -14144
rect 20120 -14177 20136 -14160
rect 19674 -14194 19876 -14177
rect 18916 -14232 19876 -14194
rect 19934 -14194 20136 -14177
rect 20692 -14177 20708 -14160
rect 21138 -14160 21726 -14144
rect 21138 -14177 21154 -14160
rect 20692 -14194 20894 -14177
rect 19934 -14232 20894 -14194
rect 20952 -14194 21154 -14177
rect 21710 -14177 21726 -14160
rect 22156 -14160 22744 -14144
rect 22156 -14177 22172 -14160
rect 21710 -14194 21912 -14177
rect 20952 -14232 21912 -14194
rect 21970 -14194 22172 -14177
rect 22728 -14177 22744 -14160
rect 22728 -14194 22930 -14177
rect 21970 -14232 22930 -14194
rect -9138 -14786 -8178 -14748
rect -9138 -14803 -8936 -14786
rect -8952 -14820 -8936 -14803
rect -8380 -14803 -8178 -14786
rect -8120 -14786 -7160 -14748
rect -8120 -14803 -7918 -14786
rect -8380 -14820 -8364 -14803
rect -8952 -14836 -8364 -14820
rect -7934 -14820 -7918 -14803
rect -7362 -14803 -7160 -14786
rect -7102 -14786 -6142 -14748
rect -7102 -14803 -6900 -14786
rect -7362 -14820 -7346 -14803
rect -7934 -14836 -7346 -14820
rect -6916 -14820 -6900 -14803
rect -6344 -14803 -6142 -14786
rect -6084 -14786 -5124 -14748
rect -6084 -14803 -5882 -14786
rect -6344 -14820 -6328 -14803
rect -6916 -14836 -6328 -14820
rect -5898 -14820 -5882 -14803
rect -5326 -14803 -5124 -14786
rect -5066 -14786 -4106 -14748
rect -5066 -14803 -4864 -14786
rect -5326 -14820 -5310 -14803
rect -5898 -14836 -5310 -14820
rect -4880 -14820 -4864 -14803
rect -4308 -14803 -4106 -14786
rect -4048 -14786 -3088 -14748
rect -4048 -14803 -3846 -14786
rect -4308 -14820 -4292 -14803
rect -4880 -14836 -4292 -14820
rect -3862 -14820 -3846 -14803
rect -3290 -14803 -3088 -14786
rect -3030 -14786 -2070 -14748
rect -3030 -14803 -2828 -14786
rect -3290 -14820 -3274 -14803
rect -3862 -14836 -3274 -14820
rect -2844 -14820 -2828 -14803
rect -2272 -14803 -2070 -14786
rect -2012 -14786 -1052 -14748
rect -2012 -14803 -1810 -14786
rect -2272 -14820 -2256 -14803
rect -2844 -14836 -2256 -14820
rect -1826 -14820 -1810 -14803
rect -1254 -14803 -1052 -14786
rect -994 -14786 -34 -14748
rect -994 -14803 -792 -14786
rect -1254 -14820 -1238 -14803
rect -1826 -14836 -1238 -14820
rect -808 -14820 -792 -14803
rect -236 -14803 -34 -14786
rect -236 -14820 -220 -14803
rect -808 -14836 -220 -14820
rect 2628 -14870 3588 -14832
rect -8952 -14894 -8364 -14878
rect -8952 -14911 -8936 -14894
rect -9138 -14928 -8936 -14911
rect -8380 -14911 -8364 -14894
rect -7934 -14894 -7346 -14878
rect -7934 -14911 -7918 -14894
rect -8380 -14928 -8178 -14911
rect -9138 -14966 -8178 -14928
rect -8120 -14928 -7918 -14911
rect -7362 -14911 -7346 -14894
rect -6916 -14894 -6328 -14878
rect -6916 -14911 -6900 -14894
rect -7362 -14928 -7160 -14911
rect -8120 -14966 -7160 -14928
rect -7102 -14928 -6900 -14911
rect -6344 -14911 -6328 -14894
rect -5898 -14894 -5310 -14878
rect -5898 -14911 -5882 -14894
rect -6344 -14928 -6142 -14911
rect -7102 -14966 -6142 -14928
rect -6084 -14928 -5882 -14911
rect -5326 -14911 -5310 -14894
rect -4880 -14894 -4292 -14878
rect -4880 -14911 -4864 -14894
rect -5326 -14928 -5124 -14911
rect -6084 -14966 -5124 -14928
rect -5066 -14928 -4864 -14911
rect -4308 -14911 -4292 -14894
rect -3862 -14894 -3274 -14878
rect -3862 -14911 -3846 -14894
rect -4308 -14928 -4106 -14911
rect -5066 -14966 -4106 -14928
rect -4048 -14928 -3846 -14911
rect -3290 -14911 -3274 -14894
rect -2844 -14894 -2256 -14878
rect -2844 -14911 -2828 -14894
rect -3290 -14928 -3088 -14911
rect -4048 -14966 -3088 -14928
rect -3030 -14928 -2828 -14911
rect -2272 -14911 -2256 -14894
rect -1826 -14894 -1238 -14878
rect -1826 -14911 -1810 -14894
rect -2272 -14928 -2070 -14911
rect -3030 -14966 -2070 -14928
rect -2012 -14928 -1810 -14911
rect -1254 -14911 -1238 -14894
rect -808 -14894 -220 -14878
rect 2628 -14887 2830 -14870
rect -808 -14911 -792 -14894
rect -1254 -14928 -1052 -14911
rect -2012 -14966 -1052 -14928
rect -994 -14928 -792 -14911
rect -236 -14911 -220 -14894
rect 2814 -14904 2830 -14887
rect 3386 -14887 3588 -14870
rect 3646 -14870 4606 -14832
rect 3646 -14887 3848 -14870
rect 3386 -14904 3402 -14887
rect -236 -14928 -34 -14911
rect 2814 -14920 3402 -14904
rect 3832 -14904 3848 -14887
rect 4404 -14887 4606 -14870
rect 4664 -14870 5624 -14832
rect 4664 -14887 4866 -14870
rect 4404 -14904 4420 -14887
rect 3832 -14920 4420 -14904
rect 4850 -14904 4866 -14887
rect 5422 -14887 5624 -14870
rect 5682 -14870 6642 -14832
rect 5682 -14887 5884 -14870
rect 5422 -14904 5438 -14887
rect 4850 -14920 5438 -14904
rect 5868 -14904 5884 -14887
rect 6440 -14887 6642 -14870
rect 6700 -14870 7660 -14832
rect 6700 -14887 6902 -14870
rect 6440 -14904 6456 -14887
rect 5868 -14920 6456 -14904
rect 6886 -14904 6902 -14887
rect 7458 -14887 7660 -14870
rect 7718 -14870 8678 -14832
rect 7718 -14887 7920 -14870
rect 7458 -14904 7474 -14887
rect 6886 -14920 7474 -14904
rect 7904 -14904 7920 -14887
rect 8476 -14887 8678 -14870
rect 8736 -14870 9696 -14832
rect 8736 -14887 8938 -14870
rect 8476 -14904 8492 -14887
rect 7904 -14920 8492 -14904
rect 8922 -14904 8938 -14887
rect 9494 -14887 9696 -14870
rect 9754 -14870 10714 -14832
rect 9754 -14887 9956 -14870
rect 9494 -14904 9510 -14887
rect 8922 -14920 9510 -14904
rect 9940 -14904 9956 -14887
rect 10512 -14887 10714 -14870
rect 10772 -14870 11732 -14832
rect 10772 -14887 10974 -14870
rect 10512 -14904 10528 -14887
rect 9940 -14920 10528 -14904
rect 10958 -14904 10974 -14887
rect 11530 -14887 11732 -14870
rect 11790 -14870 12750 -14832
rect 11790 -14887 11992 -14870
rect 11530 -14904 11546 -14887
rect 10958 -14920 11546 -14904
rect 11976 -14904 11992 -14887
rect 12548 -14887 12750 -14870
rect 12808 -14870 13768 -14832
rect 12808 -14887 13010 -14870
rect 12548 -14904 12564 -14887
rect 11976 -14920 12564 -14904
rect 12994 -14904 13010 -14887
rect 13566 -14887 13768 -14870
rect 13826 -14870 14786 -14832
rect 13826 -14887 14028 -14870
rect 13566 -14904 13582 -14887
rect 12994 -14920 13582 -14904
rect 14012 -14904 14028 -14887
rect 14584 -14887 14786 -14870
rect 14844 -14870 15804 -14832
rect 14844 -14887 15046 -14870
rect 14584 -14904 14600 -14887
rect 14012 -14920 14600 -14904
rect 15030 -14904 15046 -14887
rect 15602 -14887 15804 -14870
rect 15862 -14870 16822 -14832
rect 15862 -14887 16064 -14870
rect 15602 -14904 15618 -14887
rect 15030 -14920 15618 -14904
rect 16048 -14904 16064 -14887
rect 16620 -14887 16822 -14870
rect 16880 -14870 17840 -14832
rect 16880 -14887 17082 -14870
rect 16620 -14904 16636 -14887
rect 16048 -14920 16636 -14904
rect 17066 -14904 17082 -14887
rect 17638 -14887 17840 -14870
rect 17898 -14870 18858 -14832
rect 17898 -14887 18100 -14870
rect 17638 -14904 17654 -14887
rect 17066 -14920 17654 -14904
rect 18084 -14904 18100 -14887
rect 18656 -14887 18858 -14870
rect 18916 -14870 19876 -14832
rect 18916 -14887 19118 -14870
rect 18656 -14904 18672 -14887
rect 18084 -14920 18672 -14904
rect 19102 -14904 19118 -14887
rect 19674 -14887 19876 -14870
rect 19934 -14870 20894 -14832
rect 19934 -14887 20136 -14870
rect 19674 -14904 19690 -14887
rect 19102 -14920 19690 -14904
rect 20120 -14904 20136 -14887
rect 20692 -14887 20894 -14870
rect 20952 -14870 21912 -14832
rect 20952 -14887 21154 -14870
rect 20692 -14904 20708 -14887
rect 20120 -14920 20708 -14904
rect 21138 -14904 21154 -14887
rect 21710 -14887 21912 -14870
rect 21970 -14870 22930 -14832
rect 21970 -14887 22172 -14870
rect 21710 -14904 21726 -14887
rect 21138 -14920 21726 -14904
rect 22156 -14904 22172 -14887
rect 22728 -14887 22930 -14870
rect 22728 -14904 22744 -14887
rect 22156 -14920 22744 -14904
rect -994 -14966 -34 -14928
rect 2814 -15392 3402 -15376
rect 2814 -15409 2830 -15392
rect 2628 -15426 2830 -15409
rect 3386 -15409 3402 -15392
rect 3832 -15392 4420 -15376
rect 3832 -15409 3848 -15392
rect 3386 -15426 3588 -15409
rect 2628 -15464 3588 -15426
rect 3646 -15426 3848 -15409
rect 4404 -15409 4420 -15392
rect 4850 -15392 5438 -15376
rect 4850 -15409 4866 -15392
rect 4404 -15426 4606 -15409
rect 3646 -15464 4606 -15426
rect 4664 -15426 4866 -15409
rect 5422 -15409 5438 -15392
rect 5868 -15392 6456 -15376
rect 5868 -15409 5884 -15392
rect 5422 -15426 5624 -15409
rect 4664 -15464 5624 -15426
rect 5682 -15426 5884 -15409
rect 6440 -15409 6456 -15392
rect 6886 -15392 7474 -15376
rect 6886 -15409 6902 -15392
rect 6440 -15426 6642 -15409
rect 5682 -15464 6642 -15426
rect 6700 -15426 6902 -15409
rect 7458 -15409 7474 -15392
rect 7904 -15392 8492 -15376
rect 7904 -15409 7920 -15392
rect 7458 -15426 7660 -15409
rect 6700 -15464 7660 -15426
rect 7718 -15426 7920 -15409
rect 8476 -15409 8492 -15392
rect 8922 -15392 9510 -15376
rect 8922 -15409 8938 -15392
rect 8476 -15426 8678 -15409
rect 7718 -15464 8678 -15426
rect 8736 -15426 8938 -15409
rect 9494 -15409 9510 -15392
rect 9940 -15392 10528 -15376
rect 9940 -15409 9956 -15392
rect 9494 -15426 9696 -15409
rect 8736 -15464 9696 -15426
rect 9754 -15426 9956 -15409
rect 10512 -15409 10528 -15392
rect 10958 -15392 11546 -15376
rect 10958 -15409 10974 -15392
rect 10512 -15426 10714 -15409
rect 9754 -15464 10714 -15426
rect 10772 -15426 10974 -15409
rect 11530 -15409 11546 -15392
rect 11976 -15392 12564 -15376
rect 11976 -15409 11992 -15392
rect 11530 -15426 11732 -15409
rect 10772 -15464 11732 -15426
rect 11790 -15426 11992 -15409
rect 12548 -15409 12564 -15392
rect 12994 -15392 13582 -15376
rect 12994 -15409 13010 -15392
rect 12548 -15426 12750 -15409
rect 11790 -15464 12750 -15426
rect 12808 -15426 13010 -15409
rect 13566 -15409 13582 -15392
rect 14012 -15392 14600 -15376
rect 14012 -15409 14028 -15392
rect 13566 -15426 13768 -15409
rect 12808 -15464 13768 -15426
rect 13826 -15426 14028 -15409
rect 14584 -15409 14600 -15392
rect 15030 -15392 15618 -15376
rect 15030 -15409 15046 -15392
rect 14584 -15426 14786 -15409
rect 13826 -15464 14786 -15426
rect 14844 -15426 15046 -15409
rect 15602 -15409 15618 -15392
rect 16048 -15392 16636 -15376
rect 16048 -15409 16064 -15392
rect 15602 -15426 15804 -15409
rect 14844 -15464 15804 -15426
rect 15862 -15426 16064 -15409
rect 16620 -15409 16636 -15392
rect 17066 -15392 17654 -15376
rect 17066 -15409 17082 -15392
rect 16620 -15426 16822 -15409
rect 15862 -15464 16822 -15426
rect 16880 -15426 17082 -15409
rect 17638 -15409 17654 -15392
rect 18084 -15392 18672 -15376
rect 18084 -15409 18100 -15392
rect 17638 -15426 17840 -15409
rect 16880 -15464 17840 -15426
rect 17898 -15426 18100 -15409
rect 18656 -15409 18672 -15392
rect 19102 -15392 19690 -15376
rect 19102 -15409 19118 -15392
rect 18656 -15426 18858 -15409
rect 17898 -15464 18858 -15426
rect 18916 -15426 19118 -15409
rect 19674 -15409 19690 -15392
rect 20120 -15392 20708 -15376
rect 20120 -15409 20136 -15392
rect 19674 -15426 19876 -15409
rect 18916 -15464 19876 -15426
rect 19934 -15426 20136 -15409
rect 20692 -15409 20708 -15392
rect 21138 -15392 21726 -15376
rect 21138 -15409 21154 -15392
rect 20692 -15426 20894 -15409
rect 19934 -15464 20894 -15426
rect 20952 -15426 21154 -15409
rect 21710 -15409 21726 -15392
rect 22156 -15392 22744 -15376
rect 22156 -15409 22172 -15392
rect 21710 -15426 21912 -15409
rect 20952 -15464 21912 -15426
rect 21970 -15426 22172 -15409
rect 22728 -15409 22744 -15392
rect 22728 -15426 22930 -15409
rect 21970 -15464 22930 -15426
rect -9138 -15604 -8178 -15566
rect -9138 -15621 -8936 -15604
rect -8952 -15638 -8936 -15621
rect -8380 -15621 -8178 -15604
rect -8120 -15604 -7160 -15566
rect -8120 -15621 -7918 -15604
rect -8380 -15638 -8364 -15621
rect -8952 -15654 -8364 -15638
rect -7934 -15638 -7918 -15621
rect -7362 -15621 -7160 -15604
rect -7102 -15604 -6142 -15566
rect -7102 -15621 -6900 -15604
rect -7362 -15638 -7346 -15621
rect -7934 -15654 -7346 -15638
rect -6916 -15638 -6900 -15621
rect -6344 -15621 -6142 -15604
rect -6084 -15604 -5124 -15566
rect -6084 -15621 -5882 -15604
rect -6344 -15638 -6328 -15621
rect -6916 -15654 -6328 -15638
rect -5898 -15638 -5882 -15621
rect -5326 -15621 -5124 -15604
rect -5066 -15604 -4106 -15566
rect -5066 -15621 -4864 -15604
rect -5326 -15638 -5310 -15621
rect -5898 -15654 -5310 -15638
rect -4880 -15638 -4864 -15621
rect -4308 -15621 -4106 -15604
rect -4048 -15604 -3088 -15566
rect -4048 -15621 -3846 -15604
rect -4308 -15638 -4292 -15621
rect -4880 -15654 -4292 -15638
rect -3862 -15638 -3846 -15621
rect -3290 -15621 -3088 -15604
rect -3030 -15604 -2070 -15566
rect -3030 -15621 -2828 -15604
rect -3290 -15638 -3274 -15621
rect -3862 -15654 -3274 -15638
rect -2844 -15638 -2828 -15621
rect -2272 -15621 -2070 -15604
rect -2012 -15604 -1052 -15566
rect -2012 -15621 -1810 -15604
rect -2272 -15638 -2256 -15621
rect -2844 -15654 -2256 -15638
rect -1826 -15638 -1810 -15621
rect -1254 -15621 -1052 -15604
rect -994 -15604 -34 -15566
rect -994 -15621 -792 -15604
rect -1254 -15638 -1238 -15621
rect -1826 -15654 -1238 -15638
rect -808 -15638 -792 -15621
rect -236 -15621 -34 -15604
rect -236 -15638 -220 -15621
rect -808 -15654 -220 -15638
rect -8952 -15712 -8364 -15696
rect -8952 -15729 -8936 -15712
rect -9138 -15746 -8936 -15729
rect -8380 -15729 -8364 -15712
rect -7934 -15712 -7346 -15696
rect -7934 -15729 -7918 -15712
rect -8380 -15746 -8178 -15729
rect -9138 -15784 -8178 -15746
rect -8120 -15746 -7918 -15729
rect -7362 -15729 -7346 -15712
rect -6916 -15712 -6328 -15696
rect -6916 -15729 -6900 -15712
rect -7362 -15746 -7160 -15729
rect -8120 -15784 -7160 -15746
rect -7102 -15746 -6900 -15729
rect -6344 -15729 -6328 -15712
rect -5898 -15712 -5310 -15696
rect -5898 -15729 -5882 -15712
rect -6344 -15746 -6142 -15729
rect -7102 -15784 -6142 -15746
rect -6084 -15746 -5882 -15729
rect -5326 -15729 -5310 -15712
rect -4880 -15712 -4292 -15696
rect -4880 -15729 -4864 -15712
rect -5326 -15746 -5124 -15729
rect -6084 -15784 -5124 -15746
rect -5066 -15746 -4864 -15729
rect -4308 -15729 -4292 -15712
rect -3862 -15712 -3274 -15696
rect -3862 -15729 -3846 -15712
rect -4308 -15746 -4106 -15729
rect -5066 -15784 -4106 -15746
rect -4048 -15746 -3846 -15729
rect -3290 -15729 -3274 -15712
rect -2844 -15712 -2256 -15696
rect -2844 -15729 -2828 -15712
rect -3290 -15746 -3088 -15729
rect -4048 -15784 -3088 -15746
rect -3030 -15746 -2828 -15729
rect -2272 -15729 -2256 -15712
rect -1826 -15712 -1238 -15696
rect -1826 -15729 -1810 -15712
rect -2272 -15746 -2070 -15729
rect -3030 -15784 -2070 -15746
rect -2012 -15746 -1810 -15729
rect -1254 -15729 -1238 -15712
rect -808 -15712 -220 -15696
rect -808 -15729 -792 -15712
rect -1254 -15746 -1052 -15729
rect -2012 -15784 -1052 -15746
rect -994 -15746 -792 -15729
rect -236 -15729 -220 -15712
rect -236 -15746 -34 -15729
rect -994 -15784 -34 -15746
rect 2628 -16102 3588 -16064
rect 2628 -16119 2830 -16102
rect 2814 -16136 2830 -16119
rect 3386 -16119 3588 -16102
rect 3646 -16102 4606 -16064
rect 3646 -16119 3848 -16102
rect 3386 -16136 3402 -16119
rect 2814 -16152 3402 -16136
rect 3832 -16136 3848 -16119
rect 4404 -16119 4606 -16102
rect 4664 -16102 5624 -16064
rect 4664 -16119 4866 -16102
rect 4404 -16136 4420 -16119
rect 3832 -16152 4420 -16136
rect 4850 -16136 4866 -16119
rect 5422 -16119 5624 -16102
rect 5682 -16102 6642 -16064
rect 5682 -16119 5884 -16102
rect 5422 -16136 5438 -16119
rect 4850 -16152 5438 -16136
rect 5868 -16136 5884 -16119
rect 6440 -16119 6642 -16102
rect 6700 -16102 7660 -16064
rect 6700 -16119 6902 -16102
rect 6440 -16136 6456 -16119
rect 5868 -16152 6456 -16136
rect 6886 -16136 6902 -16119
rect 7458 -16119 7660 -16102
rect 7718 -16102 8678 -16064
rect 7718 -16119 7920 -16102
rect 7458 -16136 7474 -16119
rect 6886 -16152 7474 -16136
rect 7904 -16136 7920 -16119
rect 8476 -16119 8678 -16102
rect 8736 -16102 9696 -16064
rect 8736 -16119 8938 -16102
rect 8476 -16136 8492 -16119
rect 7904 -16152 8492 -16136
rect 8922 -16136 8938 -16119
rect 9494 -16119 9696 -16102
rect 9754 -16102 10714 -16064
rect 9754 -16119 9956 -16102
rect 9494 -16136 9510 -16119
rect 8922 -16152 9510 -16136
rect 9940 -16136 9956 -16119
rect 10512 -16119 10714 -16102
rect 10772 -16102 11732 -16064
rect 10772 -16119 10974 -16102
rect 10512 -16136 10528 -16119
rect 9940 -16152 10528 -16136
rect 10958 -16136 10974 -16119
rect 11530 -16119 11732 -16102
rect 11790 -16102 12750 -16064
rect 11790 -16119 11992 -16102
rect 11530 -16136 11546 -16119
rect 10958 -16152 11546 -16136
rect 11976 -16136 11992 -16119
rect 12548 -16119 12750 -16102
rect 12808 -16102 13768 -16064
rect 12808 -16119 13010 -16102
rect 12548 -16136 12564 -16119
rect 11976 -16152 12564 -16136
rect 12994 -16136 13010 -16119
rect 13566 -16119 13768 -16102
rect 13826 -16102 14786 -16064
rect 13826 -16119 14028 -16102
rect 13566 -16136 13582 -16119
rect 12994 -16152 13582 -16136
rect 14012 -16136 14028 -16119
rect 14584 -16119 14786 -16102
rect 14844 -16102 15804 -16064
rect 14844 -16119 15046 -16102
rect 14584 -16136 14600 -16119
rect 14012 -16152 14600 -16136
rect 15030 -16136 15046 -16119
rect 15602 -16119 15804 -16102
rect 15862 -16102 16822 -16064
rect 15862 -16119 16064 -16102
rect 15602 -16136 15618 -16119
rect 15030 -16152 15618 -16136
rect 16048 -16136 16064 -16119
rect 16620 -16119 16822 -16102
rect 16880 -16102 17840 -16064
rect 16880 -16119 17082 -16102
rect 16620 -16136 16636 -16119
rect 16048 -16152 16636 -16136
rect 17066 -16136 17082 -16119
rect 17638 -16119 17840 -16102
rect 17898 -16102 18858 -16064
rect 17898 -16119 18100 -16102
rect 17638 -16136 17654 -16119
rect 17066 -16152 17654 -16136
rect 18084 -16136 18100 -16119
rect 18656 -16119 18858 -16102
rect 18916 -16102 19876 -16064
rect 18916 -16119 19118 -16102
rect 18656 -16136 18672 -16119
rect 18084 -16152 18672 -16136
rect 19102 -16136 19118 -16119
rect 19674 -16119 19876 -16102
rect 19934 -16102 20894 -16064
rect 19934 -16119 20136 -16102
rect 19674 -16136 19690 -16119
rect 19102 -16152 19690 -16136
rect 20120 -16136 20136 -16119
rect 20692 -16119 20894 -16102
rect 20952 -16102 21912 -16064
rect 20952 -16119 21154 -16102
rect 20692 -16136 20708 -16119
rect 20120 -16152 20708 -16136
rect 21138 -16136 21154 -16119
rect 21710 -16119 21912 -16102
rect 21970 -16102 22930 -16064
rect 21970 -16119 22172 -16102
rect 21710 -16136 21726 -16119
rect 21138 -16152 21726 -16136
rect 22156 -16136 22172 -16119
rect 22728 -16119 22930 -16102
rect 22728 -16136 22744 -16119
rect 22156 -16152 22744 -16136
rect -9138 -16422 -8178 -16384
rect -9138 -16439 -8936 -16422
rect -8952 -16456 -8936 -16439
rect -8380 -16439 -8178 -16422
rect -8120 -16422 -7160 -16384
rect -8120 -16439 -7918 -16422
rect -8380 -16456 -8364 -16439
rect -8952 -16472 -8364 -16456
rect -7934 -16456 -7918 -16439
rect -7362 -16439 -7160 -16422
rect -7102 -16422 -6142 -16384
rect -7102 -16439 -6900 -16422
rect -7362 -16456 -7346 -16439
rect -7934 -16472 -7346 -16456
rect -6916 -16456 -6900 -16439
rect -6344 -16439 -6142 -16422
rect -6084 -16422 -5124 -16384
rect -6084 -16439 -5882 -16422
rect -6344 -16456 -6328 -16439
rect -6916 -16472 -6328 -16456
rect -5898 -16456 -5882 -16439
rect -5326 -16439 -5124 -16422
rect -5066 -16422 -4106 -16384
rect -5066 -16439 -4864 -16422
rect -5326 -16456 -5310 -16439
rect -5898 -16472 -5310 -16456
rect -4880 -16456 -4864 -16439
rect -4308 -16439 -4106 -16422
rect -4048 -16422 -3088 -16384
rect -4048 -16439 -3846 -16422
rect -4308 -16456 -4292 -16439
rect -4880 -16472 -4292 -16456
rect -3862 -16456 -3846 -16439
rect -3290 -16439 -3088 -16422
rect -3030 -16422 -2070 -16384
rect -3030 -16439 -2828 -16422
rect -3290 -16456 -3274 -16439
rect -3862 -16472 -3274 -16456
rect -2844 -16456 -2828 -16439
rect -2272 -16439 -2070 -16422
rect -2012 -16422 -1052 -16384
rect -2012 -16439 -1810 -16422
rect -2272 -16456 -2256 -16439
rect -2844 -16472 -2256 -16456
rect -1826 -16456 -1810 -16439
rect -1254 -16439 -1052 -16422
rect -994 -16422 -34 -16384
rect -994 -16439 -792 -16422
rect -1254 -16456 -1238 -16439
rect -1826 -16472 -1238 -16456
rect -808 -16456 -792 -16439
rect -236 -16439 -34 -16422
rect -236 -16456 -220 -16439
rect -808 -16472 -220 -16456
rect -8952 -16530 -8364 -16514
rect -8952 -16547 -8936 -16530
rect -9138 -16564 -8936 -16547
rect -8380 -16547 -8364 -16530
rect -7934 -16530 -7346 -16514
rect -7934 -16547 -7918 -16530
rect -8380 -16564 -8178 -16547
rect -9138 -16602 -8178 -16564
rect -8120 -16564 -7918 -16547
rect -7362 -16547 -7346 -16530
rect -6916 -16530 -6328 -16514
rect -6916 -16547 -6900 -16530
rect -7362 -16564 -7160 -16547
rect -8120 -16602 -7160 -16564
rect -7102 -16564 -6900 -16547
rect -6344 -16547 -6328 -16530
rect -5898 -16530 -5310 -16514
rect -5898 -16547 -5882 -16530
rect -6344 -16564 -6142 -16547
rect -7102 -16602 -6142 -16564
rect -6084 -16564 -5882 -16547
rect -5326 -16547 -5310 -16530
rect -4880 -16530 -4292 -16514
rect -4880 -16547 -4864 -16530
rect -5326 -16564 -5124 -16547
rect -6084 -16602 -5124 -16564
rect -5066 -16564 -4864 -16547
rect -4308 -16547 -4292 -16530
rect -3862 -16530 -3274 -16514
rect -3862 -16547 -3846 -16530
rect -4308 -16564 -4106 -16547
rect -5066 -16602 -4106 -16564
rect -4048 -16564 -3846 -16547
rect -3290 -16547 -3274 -16530
rect -2844 -16530 -2256 -16514
rect -2844 -16547 -2828 -16530
rect -3290 -16564 -3088 -16547
rect -4048 -16602 -3088 -16564
rect -3030 -16564 -2828 -16547
rect -2272 -16547 -2256 -16530
rect -1826 -16530 -1238 -16514
rect -1826 -16547 -1810 -16530
rect -2272 -16564 -2070 -16547
rect -3030 -16602 -2070 -16564
rect -2012 -16564 -1810 -16547
rect -1254 -16547 -1238 -16530
rect -808 -16530 -220 -16514
rect -808 -16547 -792 -16530
rect -1254 -16564 -1052 -16547
rect -2012 -16602 -1052 -16564
rect -994 -16564 -792 -16547
rect -236 -16547 -220 -16530
rect -236 -16564 -34 -16547
rect -994 -16602 -34 -16564
rect 2812 -16626 3400 -16610
rect 2812 -16643 2828 -16626
rect 2626 -16660 2828 -16643
rect 3384 -16643 3400 -16626
rect 3830 -16626 4418 -16610
rect 3830 -16643 3846 -16626
rect 3384 -16660 3586 -16643
rect 2626 -16698 3586 -16660
rect 3644 -16660 3846 -16643
rect 4402 -16643 4418 -16626
rect 4848 -16626 5436 -16610
rect 4848 -16643 4864 -16626
rect 4402 -16660 4604 -16643
rect 3644 -16698 4604 -16660
rect 4662 -16660 4864 -16643
rect 5420 -16643 5436 -16626
rect 5866 -16626 6454 -16610
rect 5866 -16643 5882 -16626
rect 5420 -16660 5622 -16643
rect 4662 -16698 5622 -16660
rect 5680 -16660 5882 -16643
rect 6438 -16643 6454 -16626
rect 6884 -16626 7472 -16610
rect 6884 -16643 6900 -16626
rect 6438 -16660 6640 -16643
rect 5680 -16698 6640 -16660
rect 6698 -16660 6900 -16643
rect 7456 -16643 7472 -16626
rect 7902 -16626 8490 -16610
rect 7902 -16643 7918 -16626
rect 7456 -16660 7658 -16643
rect 6698 -16698 7658 -16660
rect 7716 -16660 7918 -16643
rect 8474 -16643 8490 -16626
rect 8920 -16626 9508 -16610
rect 8920 -16643 8936 -16626
rect 8474 -16660 8676 -16643
rect 7716 -16698 8676 -16660
rect 8734 -16660 8936 -16643
rect 9492 -16643 9508 -16626
rect 9938 -16626 10526 -16610
rect 9938 -16643 9954 -16626
rect 9492 -16660 9694 -16643
rect 8734 -16698 9694 -16660
rect 9752 -16660 9954 -16643
rect 10510 -16643 10526 -16626
rect 10956 -16626 11544 -16610
rect 10956 -16643 10972 -16626
rect 10510 -16660 10712 -16643
rect 9752 -16698 10712 -16660
rect 10770 -16660 10972 -16643
rect 11528 -16643 11544 -16626
rect 11974 -16626 12562 -16610
rect 11974 -16643 11990 -16626
rect 11528 -16660 11730 -16643
rect 10770 -16698 11730 -16660
rect 11788 -16660 11990 -16643
rect 12546 -16643 12562 -16626
rect 12992 -16626 13580 -16610
rect 12992 -16643 13008 -16626
rect 12546 -16660 12748 -16643
rect 11788 -16698 12748 -16660
rect 12806 -16660 13008 -16643
rect 13564 -16643 13580 -16626
rect 14010 -16626 14598 -16610
rect 14010 -16643 14026 -16626
rect 13564 -16660 13766 -16643
rect 12806 -16698 13766 -16660
rect 13824 -16660 14026 -16643
rect 14582 -16643 14598 -16626
rect 15028 -16626 15616 -16610
rect 15028 -16643 15044 -16626
rect 14582 -16660 14784 -16643
rect 13824 -16698 14784 -16660
rect 14842 -16660 15044 -16643
rect 15600 -16643 15616 -16626
rect 16046 -16626 16634 -16610
rect 16046 -16643 16062 -16626
rect 15600 -16660 15802 -16643
rect 14842 -16698 15802 -16660
rect 15860 -16660 16062 -16643
rect 16618 -16643 16634 -16626
rect 17064 -16626 17652 -16610
rect 17064 -16643 17080 -16626
rect 16618 -16660 16820 -16643
rect 15860 -16698 16820 -16660
rect 16878 -16660 17080 -16643
rect 17636 -16643 17652 -16626
rect 18082 -16626 18670 -16610
rect 18082 -16643 18098 -16626
rect 17636 -16660 17838 -16643
rect 16878 -16698 17838 -16660
rect 17896 -16660 18098 -16643
rect 18654 -16643 18670 -16626
rect 19100 -16626 19688 -16610
rect 19100 -16643 19116 -16626
rect 18654 -16660 18856 -16643
rect 17896 -16698 18856 -16660
rect 18914 -16660 19116 -16643
rect 19672 -16643 19688 -16626
rect 20118 -16626 20706 -16610
rect 20118 -16643 20134 -16626
rect 19672 -16660 19874 -16643
rect 18914 -16698 19874 -16660
rect 19932 -16660 20134 -16643
rect 20690 -16643 20706 -16626
rect 21136 -16626 21724 -16610
rect 21136 -16643 21152 -16626
rect 20690 -16660 20892 -16643
rect 19932 -16698 20892 -16660
rect 20950 -16660 21152 -16643
rect 21708 -16643 21724 -16626
rect 22154 -16626 22742 -16610
rect 22154 -16643 22170 -16626
rect 21708 -16660 21910 -16643
rect 20950 -16698 21910 -16660
rect 21968 -16660 22170 -16643
rect 22726 -16643 22742 -16626
rect 22726 -16660 22928 -16643
rect 21968 -16698 22928 -16660
rect -9138 -17240 -8178 -17202
rect -9138 -17257 -8936 -17240
rect -8952 -17274 -8936 -17257
rect -8380 -17257 -8178 -17240
rect -8120 -17240 -7160 -17202
rect -8120 -17257 -7918 -17240
rect -8380 -17274 -8364 -17257
rect -8952 -17290 -8364 -17274
rect -7934 -17274 -7918 -17257
rect -7362 -17257 -7160 -17240
rect -7102 -17240 -6142 -17202
rect -7102 -17257 -6900 -17240
rect -7362 -17274 -7346 -17257
rect -7934 -17290 -7346 -17274
rect -6916 -17274 -6900 -17257
rect -6344 -17257 -6142 -17240
rect -6084 -17240 -5124 -17202
rect -6084 -17257 -5882 -17240
rect -6344 -17274 -6328 -17257
rect -6916 -17290 -6328 -17274
rect -5898 -17274 -5882 -17257
rect -5326 -17257 -5124 -17240
rect -5066 -17240 -4106 -17202
rect -5066 -17257 -4864 -17240
rect -5326 -17274 -5310 -17257
rect -5898 -17290 -5310 -17274
rect -4880 -17274 -4864 -17257
rect -4308 -17257 -4106 -17240
rect -4048 -17240 -3088 -17202
rect -4048 -17257 -3846 -17240
rect -4308 -17274 -4292 -17257
rect -4880 -17290 -4292 -17274
rect -3862 -17274 -3846 -17257
rect -3290 -17257 -3088 -17240
rect -3030 -17240 -2070 -17202
rect -3030 -17257 -2828 -17240
rect -3290 -17274 -3274 -17257
rect -3862 -17290 -3274 -17274
rect -2844 -17274 -2828 -17257
rect -2272 -17257 -2070 -17240
rect -2012 -17240 -1052 -17202
rect -2012 -17257 -1810 -17240
rect -2272 -17274 -2256 -17257
rect -2844 -17290 -2256 -17274
rect -1826 -17274 -1810 -17257
rect -1254 -17257 -1052 -17240
rect -994 -17240 -34 -17202
rect -994 -17257 -792 -17240
rect -1254 -17274 -1238 -17257
rect -1826 -17290 -1238 -17274
rect -808 -17274 -792 -17257
rect -236 -17257 -34 -17240
rect -236 -17274 -220 -17257
rect -808 -17290 -220 -17274
rect -8952 -17348 -8364 -17332
rect -8952 -17365 -8936 -17348
rect -9138 -17382 -8936 -17365
rect -8380 -17365 -8364 -17348
rect -7934 -17348 -7346 -17332
rect -7934 -17365 -7918 -17348
rect -8380 -17382 -8178 -17365
rect -9138 -17420 -8178 -17382
rect -8120 -17382 -7918 -17365
rect -7362 -17365 -7346 -17348
rect -6916 -17348 -6328 -17332
rect -6916 -17365 -6900 -17348
rect -7362 -17382 -7160 -17365
rect -8120 -17420 -7160 -17382
rect -7102 -17382 -6900 -17365
rect -6344 -17365 -6328 -17348
rect -5898 -17348 -5310 -17332
rect -5898 -17365 -5882 -17348
rect -6344 -17382 -6142 -17365
rect -7102 -17420 -6142 -17382
rect -6084 -17382 -5882 -17365
rect -5326 -17365 -5310 -17348
rect -4880 -17348 -4292 -17332
rect -4880 -17365 -4864 -17348
rect -5326 -17382 -5124 -17365
rect -6084 -17420 -5124 -17382
rect -5066 -17382 -4864 -17365
rect -4308 -17365 -4292 -17348
rect -3862 -17348 -3274 -17332
rect -3862 -17365 -3846 -17348
rect -4308 -17382 -4106 -17365
rect -5066 -17420 -4106 -17382
rect -4048 -17382 -3846 -17365
rect -3290 -17365 -3274 -17348
rect -2844 -17348 -2256 -17332
rect -2844 -17365 -2828 -17348
rect -3290 -17382 -3088 -17365
rect -4048 -17420 -3088 -17382
rect -3030 -17382 -2828 -17365
rect -2272 -17365 -2256 -17348
rect -1826 -17348 -1238 -17332
rect -1826 -17365 -1810 -17348
rect -2272 -17382 -2070 -17365
rect -3030 -17420 -2070 -17382
rect -2012 -17382 -1810 -17365
rect -1254 -17365 -1238 -17348
rect -808 -17348 -220 -17332
rect -808 -17365 -792 -17348
rect -1254 -17382 -1052 -17365
rect -2012 -17420 -1052 -17382
rect -994 -17382 -792 -17365
rect -236 -17365 -220 -17348
rect 2626 -17336 3586 -17298
rect 2626 -17353 2828 -17336
rect -236 -17382 -34 -17365
rect -994 -17420 -34 -17382
rect 2812 -17370 2828 -17353
rect 3384 -17353 3586 -17336
rect 3644 -17336 4604 -17298
rect 3644 -17353 3846 -17336
rect 3384 -17370 3400 -17353
rect 2812 -17386 3400 -17370
rect 3830 -17370 3846 -17353
rect 4402 -17353 4604 -17336
rect 4662 -17336 5622 -17298
rect 4662 -17353 4864 -17336
rect 4402 -17370 4418 -17353
rect 3830 -17386 4418 -17370
rect 4848 -17370 4864 -17353
rect 5420 -17353 5622 -17336
rect 5680 -17336 6640 -17298
rect 5680 -17353 5882 -17336
rect 5420 -17370 5436 -17353
rect 4848 -17386 5436 -17370
rect 5866 -17370 5882 -17353
rect 6438 -17353 6640 -17336
rect 6698 -17336 7658 -17298
rect 6698 -17353 6900 -17336
rect 6438 -17370 6454 -17353
rect 5866 -17386 6454 -17370
rect 6884 -17370 6900 -17353
rect 7456 -17353 7658 -17336
rect 7716 -17336 8676 -17298
rect 7716 -17353 7918 -17336
rect 7456 -17370 7472 -17353
rect 6884 -17386 7472 -17370
rect 7902 -17370 7918 -17353
rect 8474 -17353 8676 -17336
rect 8734 -17336 9694 -17298
rect 8734 -17353 8936 -17336
rect 8474 -17370 8490 -17353
rect 7902 -17386 8490 -17370
rect 8920 -17370 8936 -17353
rect 9492 -17353 9694 -17336
rect 9752 -17336 10712 -17298
rect 9752 -17353 9954 -17336
rect 9492 -17370 9508 -17353
rect 8920 -17386 9508 -17370
rect 9938 -17370 9954 -17353
rect 10510 -17353 10712 -17336
rect 10770 -17336 11730 -17298
rect 10770 -17353 10972 -17336
rect 10510 -17370 10526 -17353
rect 9938 -17386 10526 -17370
rect 10956 -17370 10972 -17353
rect 11528 -17353 11730 -17336
rect 11788 -17336 12748 -17298
rect 11788 -17353 11990 -17336
rect 11528 -17370 11544 -17353
rect 10956 -17386 11544 -17370
rect 11974 -17370 11990 -17353
rect 12546 -17353 12748 -17336
rect 12806 -17336 13766 -17298
rect 12806 -17353 13008 -17336
rect 12546 -17370 12562 -17353
rect 11974 -17386 12562 -17370
rect 12992 -17370 13008 -17353
rect 13564 -17353 13766 -17336
rect 13824 -17336 14784 -17298
rect 13824 -17353 14026 -17336
rect 13564 -17370 13580 -17353
rect 12992 -17386 13580 -17370
rect 14010 -17370 14026 -17353
rect 14582 -17353 14784 -17336
rect 14842 -17336 15802 -17298
rect 14842 -17353 15044 -17336
rect 14582 -17370 14598 -17353
rect 14010 -17386 14598 -17370
rect 15028 -17370 15044 -17353
rect 15600 -17353 15802 -17336
rect 15860 -17336 16820 -17298
rect 15860 -17353 16062 -17336
rect 15600 -17370 15616 -17353
rect 15028 -17386 15616 -17370
rect 16046 -17370 16062 -17353
rect 16618 -17353 16820 -17336
rect 16878 -17336 17838 -17298
rect 16878 -17353 17080 -17336
rect 16618 -17370 16634 -17353
rect 16046 -17386 16634 -17370
rect 17064 -17370 17080 -17353
rect 17636 -17353 17838 -17336
rect 17896 -17336 18856 -17298
rect 17896 -17353 18098 -17336
rect 17636 -17370 17652 -17353
rect 17064 -17386 17652 -17370
rect 18082 -17370 18098 -17353
rect 18654 -17353 18856 -17336
rect 18914 -17336 19874 -17298
rect 18914 -17353 19116 -17336
rect 18654 -17370 18670 -17353
rect 18082 -17386 18670 -17370
rect 19100 -17370 19116 -17353
rect 19672 -17353 19874 -17336
rect 19932 -17336 20892 -17298
rect 19932 -17353 20134 -17336
rect 19672 -17370 19688 -17353
rect 19100 -17386 19688 -17370
rect 20118 -17370 20134 -17353
rect 20690 -17353 20892 -17336
rect 20950 -17336 21910 -17298
rect 20950 -17353 21152 -17336
rect 20690 -17370 20706 -17353
rect 20118 -17386 20706 -17370
rect 21136 -17370 21152 -17353
rect 21708 -17353 21910 -17336
rect 21968 -17336 22928 -17298
rect 21968 -17353 22170 -17336
rect 21708 -17370 21724 -17353
rect 21136 -17386 21724 -17370
rect 22154 -17370 22170 -17353
rect 22726 -17353 22928 -17336
rect 22726 -17370 22742 -17353
rect 22154 -17386 22742 -17370
rect 2812 -17860 3400 -17844
rect 2812 -17877 2828 -17860
rect 2626 -17894 2828 -17877
rect 3384 -17877 3400 -17860
rect 3830 -17860 4418 -17844
rect 3830 -17877 3846 -17860
rect 3384 -17894 3586 -17877
rect 2626 -17932 3586 -17894
rect 3644 -17894 3846 -17877
rect 4402 -17877 4418 -17860
rect 4848 -17860 5436 -17844
rect 4848 -17877 4864 -17860
rect 4402 -17894 4604 -17877
rect 3644 -17932 4604 -17894
rect 4662 -17894 4864 -17877
rect 5420 -17877 5436 -17860
rect 5866 -17860 6454 -17844
rect 5866 -17877 5882 -17860
rect 5420 -17894 5622 -17877
rect 4662 -17932 5622 -17894
rect 5680 -17894 5882 -17877
rect 6438 -17877 6454 -17860
rect 6884 -17860 7472 -17844
rect 6884 -17877 6900 -17860
rect 6438 -17894 6640 -17877
rect 5680 -17932 6640 -17894
rect 6698 -17894 6900 -17877
rect 7456 -17877 7472 -17860
rect 7902 -17860 8490 -17844
rect 7902 -17877 7918 -17860
rect 7456 -17894 7658 -17877
rect 6698 -17932 7658 -17894
rect 7716 -17894 7918 -17877
rect 8474 -17877 8490 -17860
rect 8920 -17860 9508 -17844
rect 8920 -17877 8936 -17860
rect 8474 -17894 8676 -17877
rect 7716 -17932 8676 -17894
rect 8734 -17894 8936 -17877
rect 9492 -17877 9508 -17860
rect 9938 -17860 10526 -17844
rect 9938 -17877 9954 -17860
rect 9492 -17894 9694 -17877
rect 8734 -17932 9694 -17894
rect 9752 -17894 9954 -17877
rect 10510 -17877 10526 -17860
rect 10956 -17860 11544 -17844
rect 10956 -17877 10972 -17860
rect 10510 -17894 10712 -17877
rect 9752 -17932 10712 -17894
rect 10770 -17894 10972 -17877
rect 11528 -17877 11544 -17860
rect 11974 -17860 12562 -17844
rect 11974 -17877 11990 -17860
rect 11528 -17894 11730 -17877
rect 10770 -17932 11730 -17894
rect 11788 -17894 11990 -17877
rect 12546 -17877 12562 -17860
rect 12992 -17860 13580 -17844
rect 12992 -17877 13008 -17860
rect 12546 -17894 12748 -17877
rect 11788 -17932 12748 -17894
rect 12806 -17894 13008 -17877
rect 13564 -17877 13580 -17860
rect 14010 -17860 14598 -17844
rect 14010 -17877 14026 -17860
rect 13564 -17894 13766 -17877
rect 12806 -17932 13766 -17894
rect 13824 -17894 14026 -17877
rect 14582 -17877 14598 -17860
rect 15028 -17860 15616 -17844
rect 15028 -17877 15044 -17860
rect 14582 -17894 14784 -17877
rect 13824 -17932 14784 -17894
rect 14842 -17894 15044 -17877
rect 15600 -17877 15616 -17860
rect 16046 -17860 16634 -17844
rect 16046 -17877 16062 -17860
rect 15600 -17894 15802 -17877
rect 14842 -17932 15802 -17894
rect 15860 -17894 16062 -17877
rect 16618 -17877 16634 -17860
rect 17064 -17860 17652 -17844
rect 17064 -17877 17080 -17860
rect 16618 -17894 16820 -17877
rect 15860 -17932 16820 -17894
rect 16878 -17894 17080 -17877
rect 17636 -17877 17652 -17860
rect 18082 -17860 18670 -17844
rect 18082 -17877 18098 -17860
rect 17636 -17894 17838 -17877
rect 16878 -17932 17838 -17894
rect 17896 -17894 18098 -17877
rect 18654 -17877 18670 -17860
rect 19100 -17860 19688 -17844
rect 19100 -17877 19116 -17860
rect 18654 -17894 18856 -17877
rect 17896 -17932 18856 -17894
rect 18914 -17894 19116 -17877
rect 19672 -17877 19688 -17860
rect 20118 -17860 20706 -17844
rect 20118 -17877 20134 -17860
rect 19672 -17894 19874 -17877
rect 18914 -17932 19874 -17894
rect 19932 -17894 20134 -17877
rect 20690 -17877 20706 -17860
rect 21136 -17860 21724 -17844
rect 21136 -17877 21152 -17860
rect 20690 -17894 20892 -17877
rect 19932 -17932 20892 -17894
rect 20950 -17894 21152 -17877
rect 21708 -17877 21724 -17860
rect 22154 -17860 22742 -17844
rect 22154 -17877 22170 -17860
rect 21708 -17894 21910 -17877
rect 20950 -17932 21910 -17894
rect 21968 -17894 22170 -17877
rect 22726 -17877 22742 -17860
rect 22726 -17894 22928 -17877
rect 21968 -17932 22928 -17894
rect -9138 -18058 -8178 -18020
rect -9138 -18075 -8936 -18058
rect -8952 -18092 -8936 -18075
rect -8380 -18075 -8178 -18058
rect -8120 -18058 -7160 -18020
rect -8120 -18075 -7918 -18058
rect -8380 -18092 -8364 -18075
rect -8952 -18108 -8364 -18092
rect -7934 -18092 -7918 -18075
rect -7362 -18075 -7160 -18058
rect -7102 -18058 -6142 -18020
rect -7102 -18075 -6900 -18058
rect -7362 -18092 -7346 -18075
rect -7934 -18108 -7346 -18092
rect -6916 -18092 -6900 -18075
rect -6344 -18075 -6142 -18058
rect -6084 -18058 -5124 -18020
rect -6084 -18075 -5882 -18058
rect -6344 -18092 -6328 -18075
rect -6916 -18108 -6328 -18092
rect -5898 -18092 -5882 -18075
rect -5326 -18075 -5124 -18058
rect -5066 -18058 -4106 -18020
rect -5066 -18075 -4864 -18058
rect -5326 -18092 -5310 -18075
rect -5898 -18108 -5310 -18092
rect -4880 -18092 -4864 -18075
rect -4308 -18075 -4106 -18058
rect -4048 -18058 -3088 -18020
rect -4048 -18075 -3846 -18058
rect -4308 -18092 -4292 -18075
rect -4880 -18108 -4292 -18092
rect -3862 -18092 -3846 -18075
rect -3290 -18075 -3088 -18058
rect -3030 -18058 -2070 -18020
rect -3030 -18075 -2828 -18058
rect -3290 -18092 -3274 -18075
rect -3862 -18108 -3274 -18092
rect -2844 -18092 -2828 -18075
rect -2272 -18075 -2070 -18058
rect -2012 -18058 -1052 -18020
rect -2012 -18075 -1810 -18058
rect -2272 -18092 -2256 -18075
rect -2844 -18108 -2256 -18092
rect -1826 -18092 -1810 -18075
rect -1254 -18075 -1052 -18058
rect -994 -18058 -34 -18020
rect -994 -18075 -792 -18058
rect -1254 -18092 -1238 -18075
rect -1826 -18108 -1238 -18092
rect -808 -18092 -792 -18075
rect -236 -18075 -34 -18058
rect -236 -18092 -220 -18075
rect -808 -18108 -220 -18092
rect -8952 -18166 -8364 -18150
rect -8952 -18183 -8936 -18166
rect -9138 -18200 -8936 -18183
rect -8380 -18183 -8364 -18166
rect -7934 -18166 -7346 -18150
rect -7934 -18183 -7918 -18166
rect -8380 -18200 -8178 -18183
rect -9138 -18238 -8178 -18200
rect -8120 -18200 -7918 -18183
rect -7362 -18183 -7346 -18166
rect -6916 -18166 -6328 -18150
rect -6916 -18183 -6900 -18166
rect -7362 -18200 -7160 -18183
rect -8120 -18238 -7160 -18200
rect -7102 -18200 -6900 -18183
rect -6344 -18183 -6328 -18166
rect -5898 -18166 -5310 -18150
rect -5898 -18183 -5882 -18166
rect -6344 -18200 -6142 -18183
rect -7102 -18238 -6142 -18200
rect -6084 -18200 -5882 -18183
rect -5326 -18183 -5310 -18166
rect -4880 -18166 -4292 -18150
rect -4880 -18183 -4864 -18166
rect -5326 -18200 -5124 -18183
rect -6084 -18238 -5124 -18200
rect -5066 -18200 -4864 -18183
rect -4308 -18183 -4292 -18166
rect -3862 -18166 -3274 -18150
rect -3862 -18183 -3846 -18166
rect -4308 -18200 -4106 -18183
rect -5066 -18238 -4106 -18200
rect -4048 -18200 -3846 -18183
rect -3290 -18183 -3274 -18166
rect -2844 -18166 -2256 -18150
rect -2844 -18183 -2828 -18166
rect -3290 -18200 -3088 -18183
rect -4048 -18238 -3088 -18200
rect -3030 -18200 -2828 -18183
rect -2272 -18183 -2256 -18166
rect -1826 -18166 -1238 -18150
rect -1826 -18183 -1810 -18166
rect -2272 -18200 -2070 -18183
rect -3030 -18238 -2070 -18200
rect -2012 -18200 -1810 -18183
rect -1254 -18183 -1238 -18166
rect -808 -18166 -220 -18150
rect -808 -18183 -792 -18166
rect -1254 -18200 -1052 -18183
rect -2012 -18238 -1052 -18200
rect -994 -18200 -792 -18183
rect -236 -18183 -220 -18166
rect -236 -18200 -34 -18183
rect -994 -18238 -34 -18200
rect 2626 -18570 3586 -18532
rect 2626 -18587 2828 -18570
rect 2812 -18604 2828 -18587
rect 3384 -18587 3586 -18570
rect 3644 -18570 4604 -18532
rect 3644 -18587 3846 -18570
rect 3384 -18604 3400 -18587
rect 2812 -18620 3400 -18604
rect 3830 -18604 3846 -18587
rect 4402 -18587 4604 -18570
rect 4662 -18570 5622 -18532
rect 4662 -18587 4864 -18570
rect 4402 -18604 4418 -18587
rect 3830 -18620 4418 -18604
rect 4848 -18604 4864 -18587
rect 5420 -18587 5622 -18570
rect 5680 -18570 6640 -18532
rect 5680 -18587 5882 -18570
rect 5420 -18604 5436 -18587
rect 4848 -18620 5436 -18604
rect 5866 -18604 5882 -18587
rect 6438 -18587 6640 -18570
rect 6698 -18570 7658 -18532
rect 6698 -18587 6900 -18570
rect 6438 -18604 6454 -18587
rect 5866 -18620 6454 -18604
rect 6884 -18604 6900 -18587
rect 7456 -18587 7658 -18570
rect 7716 -18570 8676 -18532
rect 7716 -18587 7918 -18570
rect 7456 -18604 7472 -18587
rect 6884 -18620 7472 -18604
rect 7902 -18604 7918 -18587
rect 8474 -18587 8676 -18570
rect 8734 -18570 9694 -18532
rect 8734 -18587 8936 -18570
rect 8474 -18604 8490 -18587
rect 7902 -18620 8490 -18604
rect 8920 -18604 8936 -18587
rect 9492 -18587 9694 -18570
rect 9752 -18570 10712 -18532
rect 9752 -18587 9954 -18570
rect 9492 -18604 9508 -18587
rect 8920 -18620 9508 -18604
rect 9938 -18604 9954 -18587
rect 10510 -18587 10712 -18570
rect 10770 -18570 11730 -18532
rect 10770 -18587 10972 -18570
rect 10510 -18604 10526 -18587
rect 9938 -18620 10526 -18604
rect 10956 -18604 10972 -18587
rect 11528 -18587 11730 -18570
rect 11788 -18570 12748 -18532
rect 11788 -18587 11990 -18570
rect 11528 -18604 11544 -18587
rect 10956 -18620 11544 -18604
rect 11974 -18604 11990 -18587
rect 12546 -18587 12748 -18570
rect 12806 -18570 13766 -18532
rect 12806 -18587 13008 -18570
rect 12546 -18604 12562 -18587
rect 11974 -18620 12562 -18604
rect 12992 -18604 13008 -18587
rect 13564 -18587 13766 -18570
rect 13824 -18570 14784 -18532
rect 13824 -18587 14026 -18570
rect 13564 -18604 13580 -18587
rect 12992 -18620 13580 -18604
rect 14010 -18604 14026 -18587
rect 14582 -18587 14784 -18570
rect 14842 -18570 15802 -18532
rect 14842 -18587 15044 -18570
rect 14582 -18604 14598 -18587
rect 14010 -18620 14598 -18604
rect 15028 -18604 15044 -18587
rect 15600 -18587 15802 -18570
rect 15860 -18570 16820 -18532
rect 15860 -18587 16062 -18570
rect 15600 -18604 15616 -18587
rect 15028 -18620 15616 -18604
rect 16046 -18604 16062 -18587
rect 16618 -18587 16820 -18570
rect 16878 -18570 17838 -18532
rect 16878 -18587 17080 -18570
rect 16618 -18604 16634 -18587
rect 16046 -18620 16634 -18604
rect 17064 -18604 17080 -18587
rect 17636 -18587 17838 -18570
rect 17896 -18570 18856 -18532
rect 17896 -18587 18098 -18570
rect 17636 -18604 17652 -18587
rect 17064 -18620 17652 -18604
rect 18082 -18604 18098 -18587
rect 18654 -18587 18856 -18570
rect 18914 -18570 19874 -18532
rect 18914 -18587 19116 -18570
rect 18654 -18604 18670 -18587
rect 18082 -18620 18670 -18604
rect 19100 -18604 19116 -18587
rect 19672 -18587 19874 -18570
rect 19932 -18570 20892 -18532
rect 19932 -18587 20134 -18570
rect 19672 -18604 19688 -18587
rect 19100 -18620 19688 -18604
rect 20118 -18604 20134 -18587
rect 20690 -18587 20892 -18570
rect 20950 -18570 21910 -18532
rect 20950 -18587 21152 -18570
rect 20690 -18604 20706 -18587
rect 20118 -18620 20706 -18604
rect 21136 -18604 21152 -18587
rect 21708 -18587 21910 -18570
rect 21968 -18570 22928 -18532
rect 21968 -18587 22170 -18570
rect 21708 -18604 21724 -18587
rect 21136 -18620 21724 -18604
rect 22154 -18604 22170 -18587
rect 22726 -18587 22928 -18570
rect 22726 -18604 22742 -18587
rect 22154 -18620 22742 -18604
rect -9138 -18876 -8178 -18838
rect -9138 -18893 -8936 -18876
rect -8952 -18910 -8936 -18893
rect -8380 -18893 -8178 -18876
rect -8120 -18876 -7160 -18838
rect -8120 -18893 -7918 -18876
rect -8380 -18910 -8364 -18893
rect -8952 -18926 -8364 -18910
rect -7934 -18910 -7918 -18893
rect -7362 -18893 -7160 -18876
rect -7102 -18876 -6142 -18838
rect -7102 -18893 -6900 -18876
rect -7362 -18910 -7346 -18893
rect -7934 -18926 -7346 -18910
rect -6916 -18910 -6900 -18893
rect -6344 -18893 -6142 -18876
rect -6084 -18876 -5124 -18838
rect -6084 -18893 -5882 -18876
rect -6344 -18910 -6328 -18893
rect -6916 -18926 -6328 -18910
rect -5898 -18910 -5882 -18893
rect -5326 -18893 -5124 -18876
rect -5066 -18876 -4106 -18838
rect -5066 -18893 -4864 -18876
rect -5326 -18910 -5310 -18893
rect -5898 -18926 -5310 -18910
rect -4880 -18910 -4864 -18893
rect -4308 -18893 -4106 -18876
rect -4048 -18876 -3088 -18838
rect -4048 -18893 -3846 -18876
rect -4308 -18910 -4292 -18893
rect -4880 -18926 -4292 -18910
rect -3862 -18910 -3846 -18893
rect -3290 -18893 -3088 -18876
rect -3030 -18876 -2070 -18838
rect -3030 -18893 -2828 -18876
rect -3290 -18910 -3274 -18893
rect -3862 -18926 -3274 -18910
rect -2844 -18910 -2828 -18893
rect -2272 -18893 -2070 -18876
rect -2012 -18876 -1052 -18838
rect -2012 -18893 -1810 -18876
rect -2272 -18910 -2256 -18893
rect -2844 -18926 -2256 -18910
rect -1826 -18910 -1810 -18893
rect -1254 -18893 -1052 -18876
rect -994 -18876 -34 -18838
rect -994 -18893 -792 -18876
rect -1254 -18910 -1238 -18893
rect -1826 -18926 -1238 -18910
rect -808 -18910 -792 -18893
rect -236 -18893 -34 -18876
rect -236 -18910 -220 -18893
rect -808 -18926 -220 -18910
rect 2812 -19092 3400 -19076
rect 2812 -19109 2828 -19092
rect 2626 -19126 2828 -19109
rect 3384 -19109 3400 -19092
rect 3830 -19092 4418 -19076
rect 3830 -19109 3846 -19092
rect 3384 -19126 3586 -19109
rect 2626 -19164 3586 -19126
rect 3644 -19126 3846 -19109
rect 4402 -19109 4418 -19092
rect 4848 -19092 5436 -19076
rect 4848 -19109 4864 -19092
rect 4402 -19126 4604 -19109
rect 3644 -19164 4604 -19126
rect 4662 -19126 4864 -19109
rect 5420 -19109 5436 -19092
rect 5866 -19092 6454 -19076
rect 5866 -19109 5882 -19092
rect 5420 -19126 5622 -19109
rect 4662 -19164 5622 -19126
rect 5680 -19126 5882 -19109
rect 6438 -19109 6454 -19092
rect 6884 -19092 7472 -19076
rect 6884 -19109 6900 -19092
rect 6438 -19126 6640 -19109
rect 5680 -19164 6640 -19126
rect 6698 -19126 6900 -19109
rect 7456 -19109 7472 -19092
rect 7902 -19092 8490 -19076
rect 7902 -19109 7918 -19092
rect 7456 -19126 7658 -19109
rect 6698 -19164 7658 -19126
rect 7716 -19126 7918 -19109
rect 8474 -19109 8490 -19092
rect 8920 -19092 9508 -19076
rect 8920 -19109 8936 -19092
rect 8474 -19126 8676 -19109
rect 7716 -19164 8676 -19126
rect 8734 -19126 8936 -19109
rect 9492 -19109 9508 -19092
rect 9938 -19092 10526 -19076
rect 9938 -19109 9954 -19092
rect 9492 -19126 9694 -19109
rect 8734 -19164 9694 -19126
rect 9752 -19126 9954 -19109
rect 10510 -19109 10526 -19092
rect 10956 -19092 11544 -19076
rect 10956 -19109 10972 -19092
rect 10510 -19126 10712 -19109
rect 9752 -19164 10712 -19126
rect 10770 -19126 10972 -19109
rect 11528 -19109 11544 -19092
rect 11974 -19092 12562 -19076
rect 11974 -19109 11990 -19092
rect 11528 -19126 11730 -19109
rect 10770 -19164 11730 -19126
rect 11788 -19126 11990 -19109
rect 12546 -19109 12562 -19092
rect 12992 -19092 13580 -19076
rect 12992 -19109 13008 -19092
rect 12546 -19126 12748 -19109
rect 11788 -19164 12748 -19126
rect 12806 -19126 13008 -19109
rect 13564 -19109 13580 -19092
rect 14010 -19092 14598 -19076
rect 14010 -19109 14026 -19092
rect 13564 -19126 13766 -19109
rect 12806 -19164 13766 -19126
rect 13824 -19126 14026 -19109
rect 14582 -19109 14598 -19092
rect 15028 -19092 15616 -19076
rect 15028 -19109 15044 -19092
rect 14582 -19126 14784 -19109
rect 13824 -19164 14784 -19126
rect 14842 -19126 15044 -19109
rect 15600 -19109 15616 -19092
rect 16046 -19092 16634 -19076
rect 16046 -19109 16062 -19092
rect 15600 -19126 15802 -19109
rect 14842 -19164 15802 -19126
rect 15860 -19126 16062 -19109
rect 16618 -19109 16634 -19092
rect 17064 -19092 17652 -19076
rect 17064 -19109 17080 -19092
rect 16618 -19126 16820 -19109
rect 15860 -19164 16820 -19126
rect 16878 -19126 17080 -19109
rect 17636 -19109 17652 -19092
rect 18082 -19092 18670 -19076
rect 18082 -19109 18098 -19092
rect 17636 -19126 17838 -19109
rect 16878 -19164 17838 -19126
rect 17896 -19126 18098 -19109
rect 18654 -19109 18670 -19092
rect 19100 -19092 19688 -19076
rect 19100 -19109 19116 -19092
rect 18654 -19126 18856 -19109
rect 17896 -19164 18856 -19126
rect 18914 -19126 19116 -19109
rect 19672 -19109 19688 -19092
rect 20118 -19092 20706 -19076
rect 20118 -19109 20134 -19092
rect 19672 -19126 19874 -19109
rect 18914 -19164 19874 -19126
rect 19932 -19126 20134 -19109
rect 20690 -19109 20706 -19092
rect 21136 -19092 21724 -19076
rect 21136 -19109 21152 -19092
rect 20690 -19126 20892 -19109
rect 19932 -19164 20892 -19126
rect 20950 -19126 21152 -19109
rect 21708 -19109 21724 -19092
rect 22154 -19092 22742 -19076
rect 22154 -19109 22170 -19092
rect 21708 -19126 21910 -19109
rect 20950 -19164 21910 -19126
rect 21968 -19126 22170 -19109
rect 22726 -19109 22742 -19092
rect 22726 -19126 22928 -19109
rect 21968 -19164 22928 -19126
rect 2626 -19802 3586 -19764
rect 2626 -19819 2828 -19802
rect 2812 -19836 2828 -19819
rect 3384 -19819 3586 -19802
rect 3644 -19802 4604 -19764
rect 3644 -19819 3846 -19802
rect 3384 -19836 3400 -19819
rect 2812 -19852 3400 -19836
rect 3830 -19836 3846 -19819
rect 4402 -19819 4604 -19802
rect 4662 -19802 5622 -19764
rect 4662 -19819 4864 -19802
rect 4402 -19836 4418 -19819
rect 3830 -19852 4418 -19836
rect 4848 -19836 4864 -19819
rect 5420 -19819 5622 -19802
rect 5680 -19802 6640 -19764
rect 5680 -19819 5882 -19802
rect 5420 -19836 5436 -19819
rect 4848 -19852 5436 -19836
rect 5866 -19836 5882 -19819
rect 6438 -19819 6640 -19802
rect 6698 -19802 7658 -19764
rect 6698 -19819 6900 -19802
rect 6438 -19836 6454 -19819
rect 5866 -19852 6454 -19836
rect 6884 -19836 6900 -19819
rect 7456 -19819 7658 -19802
rect 7716 -19802 8676 -19764
rect 7716 -19819 7918 -19802
rect 7456 -19836 7472 -19819
rect 6884 -19852 7472 -19836
rect 7902 -19836 7918 -19819
rect 8474 -19819 8676 -19802
rect 8734 -19802 9694 -19764
rect 8734 -19819 8936 -19802
rect 8474 -19836 8490 -19819
rect 7902 -19852 8490 -19836
rect 8920 -19836 8936 -19819
rect 9492 -19819 9694 -19802
rect 9752 -19802 10712 -19764
rect 9752 -19819 9954 -19802
rect 9492 -19836 9508 -19819
rect 8920 -19852 9508 -19836
rect 9938 -19836 9954 -19819
rect 10510 -19819 10712 -19802
rect 10770 -19802 11730 -19764
rect 10770 -19819 10972 -19802
rect 10510 -19836 10526 -19819
rect 9938 -19852 10526 -19836
rect 10956 -19836 10972 -19819
rect 11528 -19819 11730 -19802
rect 11788 -19802 12748 -19764
rect 11788 -19819 11990 -19802
rect 11528 -19836 11544 -19819
rect 10956 -19852 11544 -19836
rect 11974 -19836 11990 -19819
rect 12546 -19819 12748 -19802
rect 12806 -19802 13766 -19764
rect 12806 -19819 13008 -19802
rect 12546 -19836 12562 -19819
rect 11974 -19852 12562 -19836
rect 12992 -19836 13008 -19819
rect 13564 -19819 13766 -19802
rect 13824 -19802 14784 -19764
rect 13824 -19819 14026 -19802
rect 13564 -19836 13580 -19819
rect 12992 -19852 13580 -19836
rect 14010 -19836 14026 -19819
rect 14582 -19819 14784 -19802
rect 14842 -19802 15802 -19764
rect 14842 -19819 15044 -19802
rect 14582 -19836 14598 -19819
rect 14010 -19852 14598 -19836
rect 15028 -19836 15044 -19819
rect 15600 -19819 15802 -19802
rect 15860 -19802 16820 -19764
rect 15860 -19819 16062 -19802
rect 15600 -19836 15616 -19819
rect 15028 -19852 15616 -19836
rect 16046 -19836 16062 -19819
rect 16618 -19819 16820 -19802
rect 16878 -19802 17838 -19764
rect 16878 -19819 17080 -19802
rect 16618 -19836 16634 -19819
rect 16046 -19852 16634 -19836
rect 17064 -19836 17080 -19819
rect 17636 -19819 17838 -19802
rect 17896 -19802 18856 -19764
rect 17896 -19819 18098 -19802
rect 17636 -19836 17652 -19819
rect 17064 -19852 17652 -19836
rect 18082 -19836 18098 -19819
rect 18654 -19819 18856 -19802
rect 18914 -19802 19874 -19764
rect 18914 -19819 19116 -19802
rect 18654 -19836 18670 -19819
rect 18082 -19852 18670 -19836
rect 19100 -19836 19116 -19819
rect 19672 -19819 19874 -19802
rect 19932 -19802 20892 -19764
rect 19932 -19819 20134 -19802
rect 19672 -19836 19688 -19819
rect 19100 -19852 19688 -19836
rect 20118 -19836 20134 -19819
rect 20690 -19819 20892 -19802
rect 20950 -19802 21910 -19764
rect 20950 -19819 21152 -19802
rect 20690 -19836 20706 -19819
rect 20118 -19852 20706 -19836
rect 21136 -19836 21152 -19819
rect 21708 -19819 21910 -19802
rect 21968 -19802 22928 -19764
rect 21968 -19819 22170 -19802
rect 21708 -19836 21724 -19819
rect 21136 -19852 21724 -19836
rect 22154 -19836 22170 -19819
rect 22726 -19819 22928 -19802
rect 22726 -19836 22742 -19819
rect 22154 -19852 22742 -19836
rect 2812 -20326 3400 -20310
rect 2812 -20343 2828 -20326
rect 2626 -20360 2828 -20343
rect 3384 -20343 3400 -20326
rect 3830 -20326 4418 -20310
rect 3830 -20343 3846 -20326
rect 3384 -20360 3586 -20343
rect 2626 -20398 3586 -20360
rect 3644 -20360 3846 -20343
rect 4402 -20343 4418 -20326
rect 4848 -20326 5436 -20310
rect 4848 -20343 4864 -20326
rect 4402 -20360 4604 -20343
rect 3644 -20398 4604 -20360
rect 4662 -20360 4864 -20343
rect 5420 -20343 5436 -20326
rect 5866 -20326 6454 -20310
rect 5866 -20343 5882 -20326
rect 5420 -20360 5622 -20343
rect 4662 -20398 5622 -20360
rect 5680 -20360 5882 -20343
rect 6438 -20343 6454 -20326
rect 6884 -20326 7472 -20310
rect 6884 -20343 6900 -20326
rect 6438 -20360 6640 -20343
rect 5680 -20398 6640 -20360
rect 6698 -20360 6900 -20343
rect 7456 -20343 7472 -20326
rect 7902 -20326 8490 -20310
rect 7902 -20343 7918 -20326
rect 7456 -20360 7658 -20343
rect 6698 -20398 7658 -20360
rect 7716 -20360 7918 -20343
rect 8474 -20343 8490 -20326
rect 8920 -20326 9508 -20310
rect 8920 -20343 8936 -20326
rect 8474 -20360 8676 -20343
rect 7716 -20398 8676 -20360
rect 8734 -20360 8936 -20343
rect 9492 -20343 9508 -20326
rect 9938 -20326 10526 -20310
rect 9938 -20343 9954 -20326
rect 9492 -20360 9694 -20343
rect 8734 -20398 9694 -20360
rect 9752 -20360 9954 -20343
rect 10510 -20343 10526 -20326
rect 10956 -20326 11544 -20310
rect 10956 -20343 10972 -20326
rect 10510 -20360 10712 -20343
rect 9752 -20398 10712 -20360
rect 10770 -20360 10972 -20343
rect 11528 -20343 11544 -20326
rect 11974 -20326 12562 -20310
rect 11974 -20343 11990 -20326
rect 11528 -20360 11730 -20343
rect 10770 -20398 11730 -20360
rect 11788 -20360 11990 -20343
rect 12546 -20343 12562 -20326
rect 12992 -20326 13580 -20310
rect 12992 -20343 13008 -20326
rect 12546 -20360 12748 -20343
rect 11788 -20398 12748 -20360
rect 12806 -20360 13008 -20343
rect 13564 -20343 13580 -20326
rect 14010 -20326 14598 -20310
rect 14010 -20343 14026 -20326
rect 13564 -20360 13766 -20343
rect 12806 -20398 13766 -20360
rect 13824 -20360 14026 -20343
rect 14582 -20343 14598 -20326
rect 15028 -20326 15616 -20310
rect 15028 -20343 15044 -20326
rect 14582 -20360 14784 -20343
rect 13824 -20398 14784 -20360
rect 14842 -20360 15044 -20343
rect 15600 -20343 15616 -20326
rect 16046 -20326 16634 -20310
rect 16046 -20343 16062 -20326
rect 15600 -20360 15802 -20343
rect 14842 -20398 15802 -20360
rect 15860 -20360 16062 -20343
rect 16618 -20343 16634 -20326
rect 17064 -20326 17652 -20310
rect 17064 -20343 17080 -20326
rect 16618 -20360 16820 -20343
rect 15860 -20398 16820 -20360
rect 16878 -20360 17080 -20343
rect 17636 -20343 17652 -20326
rect 18082 -20326 18670 -20310
rect 18082 -20343 18098 -20326
rect 17636 -20360 17838 -20343
rect 16878 -20398 17838 -20360
rect 17896 -20360 18098 -20343
rect 18654 -20343 18670 -20326
rect 19100 -20326 19688 -20310
rect 19100 -20343 19116 -20326
rect 18654 -20360 18856 -20343
rect 17896 -20398 18856 -20360
rect 18914 -20360 19116 -20343
rect 19672 -20343 19688 -20326
rect 20118 -20326 20706 -20310
rect 20118 -20343 20134 -20326
rect 19672 -20360 19874 -20343
rect 18914 -20398 19874 -20360
rect 19932 -20360 20134 -20343
rect 20690 -20343 20706 -20326
rect 21136 -20326 21724 -20310
rect 21136 -20343 21152 -20326
rect 20690 -20360 20892 -20343
rect 19932 -20398 20892 -20360
rect 20950 -20360 21152 -20343
rect 21708 -20343 21724 -20326
rect 22154 -20326 22742 -20310
rect 22154 -20343 22170 -20326
rect 21708 -20360 21910 -20343
rect 20950 -20398 21910 -20360
rect 21968 -20360 22170 -20343
rect 22726 -20343 22742 -20326
rect 22726 -20360 22928 -20343
rect 21968 -20398 22928 -20360
rect 2626 -21036 3586 -20998
rect 2626 -21053 2828 -21036
rect 2812 -21070 2828 -21053
rect 3384 -21053 3586 -21036
rect 3644 -21036 4604 -20998
rect 3644 -21053 3846 -21036
rect 3384 -21070 3400 -21053
rect 2812 -21086 3400 -21070
rect 3830 -21070 3846 -21053
rect 4402 -21053 4604 -21036
rect 4662 -21036 5622 -20998
rect 4662 -21053 4864 -21036
rect 4402 -21070 4418 -21053
rect 3830 -21086 4418 -21070
rect 4848 -21070 4864 -21053
rect 5420 -21053 5622 -21036
rect 5680 -21036 6640 -20998
rect 5680 -21053 5882 -21036
rect 5420 -21070 5436 -21053
rect 4848 -21086 5436 -21070
rect 5866 -21070 5882 -21053
rect 6438 -21053 6640 -21036
rect 6698 -21036 7658 -20998
rect 6698 -21053 6900 -21036
rect 6438 -21070 6454 -21053
rect 5866 -21086 6454 -21070
rect 6884 -21070 6900 -21053
rect 7456 -21053 7658 -21036
rect 7716 -21036 8676 -20998
rect 7716 -21053 7918 -21036
rect 7456 -21070 7472 -21053
rect 6884 -21086 7472 -21070
rect 7902 -21070 7918 -21053
rect 8474 -21053 8676 -21036
rect 8734 -21036 9694 -20998
rect 8734 -21053 8936 -21036
rect 8474 -21070 8490 -21053
rect 7902 -21086 8490 -21070
rect 8920 -21070 8936 -21053
rect 9492 -21053 9694 -21036
rect 9752 -21036 10712 -20998
rect 9752 -21053 9954 -21036
rect 9492 -21070 9508 -21053
rect 8920 -21086 9508 -21070
rect 9938 -21070 9954 -21053
rect 10510 -21053 10712 -21036
rect 10770 -21036 11730 -20998
rect 10770 -21053 10972 -21036
rect 10510 -21070 10526 -21053
rect 9938 -21086 10526 -21070
rect 10956 -21070 10972 -21053
rect 11528 -21053 11730 -21036
rect 11788 -21036 12748 -20998
rect 11788 -21053 11990 -21036
rect 11528 -21070 11544 -21053
rect 10956 -21086 11544 -21070
rect 11974 -21070 11990 -21053
rect 12546 -21053 12748 -21036
rect 12806 -21036 13766 -20998
rect 12806 -21053 13008 -21036
rect 12546 -21070 12562 -21053
rect 11974 -21086 12562 -21070
rect 12992 -21070 13008 -21053
rect 13564 -21053 13766 -21036
rect 13824 -21036 14784 -20998
rect 13824 -21053 14026 -21036
rect 13564 -21070 13580 -21053
rect 12992 -21086 13580 -21070
rect 14010 -21070 14026 -21053
rect 14582 -21053 14784 -21036
rect 14842 -21036 15802 -20998
rect 14842 -21053 15044 -21036
rect 14582 -21070 14598 -21053
rect 14010 -21086 14598 -21070
rect 15028 -21070 15044 -21053
rect 15600 -21053 15802 -21036
rect 15860 -21036 16820 -20998
rect 15860 -21053 16062 -21036
rect 15600 -21070 15616 -21053
rect 15028 -21086 15616 -21070
rect 16046 -21070 16062 -21053
rect 16618 -21053 16820 -21036
rect 16878 -21036 17838 -20998
rect 16878 -21053 17080 -21036
rect 16618 -21070 16634 -21053
rect 16046 -21086 16634 -21070
rect 17064 -21070 17080 -21053
rect 17636 -21053 17838 -21036
rect 17896 -21036 18856 -20998
rect 17896 -21053 18098 -21036
rect 17636 -21070 17652 -21053
rect 17064 -21086 17652 -21070
rect 18082 -21070 18098 -21053
rect 18654 -21053 18856 -21036
rect 18914 -21036 19874 -20998
rect 18914 -21053 19116 -21036
rect 18654 -21070 18670 -21053
rect 18082 -21086 18670 -21070
rect 19100 -21070 19116 -21053
rect 19672 -21053 19874 -21036
rect 19932 -21036 20892 -20998
rect 19932 -21053 20134 -21036
rect 19672 -21070 19688 -21053
rect 19100 -21086 19688 -21070
rect 20118 -21070 20134 -21053
rect 20690 -21053 20892 -21036
rect 20950 -21036 21910 -20998
rect 20950 -21053 21152 -21036
rect 20690 -21070 20706 -21053
rect 20118 -21086 20706 -21070
rect 21136 -21070 21152 -21053
rect 21708 -21053 21910 -21036
rect 21968 -21036 22928 -20998
rect 21968 -21053 22170 -21036
rect 21708 -21070 21724 -21053
rect 21136 -21086 21724 -21070
rect 22154 -21070 22170 -21053
rect 22726 -21053 22928 -21036
rect 22726 -21070 22742 -21053
rect 22154 -21086 22742 -21070
rect 2812 -21560 3400 -21544
rect 2812 -21577 2828 -21560
rect 2626 -21594 2828 -21577
rect 3384 -21577 3400 -21560
rect 3830 -21560 4418 -21544
rect 3830 -21577 3846 -21560
rect 3384 -21594 3586 -21577
rect 2626 -21632 3586 -21594
rect 3644 -21594 3846 -21577
rect 4402 -21577 4418 -21560
rect 4848 -21560 5436 -21544
rect 4848 -21577 4864 -21560
rect 4402 -21594 4604 -21577
rect 3644 -21632 4604 -21594
rect 4662 -21594 4864 -21577
rect 5420 -21577 5436 -21560
rect 5866 -21560 6454 -21544
rect 5866 -21577 5882 -21560
rect 5420 -21594 5622 -21577
rect 4662 -21632 5622 -21594
rect 5680 -21594 5882 -21577
rect 6438 -21577 6454 -21560
rect 6884 -21560 7472 -21544
rect 6884 -21577 6900 -21560
rect 6438 -21594 6640 -21577
rect 5680 -21632 6640 -21594
rect 6698 -21594 6900 -21577
rect 7456 -21577 7472 -21560
rect 7902 -21560 8490 -21544
rect 7902 -21577 7918 -21560
rect 7456 -21594 7658 -21577
rect 6698 -21632 7658 -21594
rect 7716 -21594 7918 -21577
rect 8474 -21577 8490 -21560
rect 8920 -21560 9508 -21544
rect 8920 -21577 8936 -21560
rect 8474 -21594 8676 -21577
rect 7716 -21632 8676 -21594
rect 8734 -21594 8936 -21577
rect 9492 -21577 9508 -21560
rect 9938 -21560 10526 -21544
rect 9938 -21577 9954 -21560
rect 9492 -21594 9694 -21577
rect 8734 -21632 9694 -21594
rect 9752 -21594 9954 -21577
rect 10510 -21577 10526 -21560
rect 10956 -21560 11544 -21544
rect 10956 -21577 10972 -21560
rect 10510 -21594 10712 -21577
rect 9752 -21632 10712 -21594
rect 10770 -21594 10972 -21577
rect 11528 -21577 11544 -21560
rect 11974 -21560 12562 -21544
rect 11974 -21577 11990 -21560
rect 11528 -21594 11730 -21577
rect 10770 -21632 11730 -21594
rect 11788 -21594 11990 -21577
rect 12546 -21577 12562 -21560
rect 12992 -21560 13580 -21544
rect 12992 -21577 13008 -21560
rect 12546 -21594 12748 -21577
rect 11788 -21632 12748 -21594
rect 12806 -21594 13008 -21577
rect 13564 -21577 13580 -21560
rect 14010 -21560 14598 -21544
rect 14010 -21577 14026 -21560
rect 13564 -21594 13766 -21577
rect 12806 -21632 13766 -21594
rect 13824 -21594 14026 -21577
rect 14582 -21577 14598 -21560
rect 15028 -21560 15616 -21544
rect 15028 -21577 15044 -21560
rect 14582 -21594 14784 -21577
rect 13824 -21632 14784 -21594
rect 14842 -21594 15044 -21577
rect 15600 -21577 15616 -21560
rect 16046 -21560 16634 -21544
rect 16046 -21577 16062 -21560
rect 15600 -21594 15802 -21577
rect 14842 -21632 15802 -21594
rect 15860 -21594 16062 -21577
rect 16618 -21577 16634 -21560
rect 17064 -21560 17652 -21544
rect 17064 -21577 17080 -21560
rect 16618 -21594 16820 -21577
rect 15860 -21632 16820 -21594
rect 16878 -21594 17080 -21577
rect 17636 -21577 17652 -21560
rect 18082 -21560 18670 -21544
rect 18082 -21577 18098 -21560
rect 17636 -21594 17838 -21577
rect 16878 -21632 17838 -21594
rect 17896 -21594 18098 -21577
rect 18654 -21577 18670 -21560
rect 19100 -21560 19688 -21544
rect 19100 -21577 19116 -21560
rect 18654 -21594 18856 -21577
rect 17896 -21632 18856 -21594
rect 18914 -21594 19116 -21577
rect 19672 -21577 19688 -21560
rect 20118 -21560 20706 -21544
rect 20118 -21577 20134 -21560
rect 19672 -21594 19874 -21577
rect 18914 -21632 19874 -21594
rect 19932 -21594 20134 -21577
rect 20690 -21577 20706 -21560
rect 21136 -21560 21724 -21544
rect 21136 -21577 21152 -21560
rect 20690 -21594 20892 -21577
rect 19932 -21632 20892 -21594
rect 20950 -21594 21152 -21577
rect 21708 -21577 21724 -21560
rect 22154 -21560 22742 -21544
rect 22154 -21577 22170 -21560
rect 21708 -21594 21910 -21577
rect 20950 -21632 21910 -21594
rect 21968 -21594 22170 -21577
rect 22726 -21577 22742 -21560
rect 22726 -21594 22928 -21577
rect 21968 -21632 22928 -21594
rect 2626 -22270 3586 -22232
rect 2626 -22287 2828 -22270
rect 2812 -22304 2828 -22287
rect 3384 -22287 3586 -22270
rect 3644 -22270 4604 -22232
rect 3644 -22287 3846 -22270
rect 3384 -22304 3400 -22287
rect 2812 -22320 3400 -22304
rect 3830 -22304 3846 -22287
rect 4402 -22287 4604 -22270
rect 4662 -22270 5622 -22232
rect 4662 -22287 4864 -22270
rect 4402 -22304 4418 -22287
rect 3830 -22320 4418 -22304
rect 4848 -22304 4864 -22287
rect 5420 -22287 5622 -22270
rect 5680 -22270 6640 -22232
rect 5680 -22287 5882 -22270
rect 5420 -22304 5436 -22287
rect 4848 -22320 5436 -22304
rect 5866 -22304 5882 -22287
rect 6438 -22287 6640 -22270
rect 6698 -22270 7658 -22232
rect 6698 -22287 6900 -22270
rect 6438 -22304 6454 -22287
rect 5866 -22320 6454 -22304
rect 6884 -22304 6900 -22287
rect 7456 -22287 7658 -22270
rect 7716 -22270 8676 -22232
rect 7716 -22287 7918 -22270
rect 7456 -22304 7472 -22287
rect 6884 -22320 7472 -22304
rect 7902 -22304 7918 -22287
rect 8474 -22287 8676 -22270
rect 8734 -22270 9694 -22232
rect 8734 -22287 8936 -22270
rect 8474 -22304 8490 -22287
rect 7902 -22320 8490 -22304
rect 8920 -22304 8936 -22287
rect 9492 -22287 9694 -22270
rect 9752 -22270 10712 -22232
rect 9752 -22287 9954 -22270
rect 9492 -22304 9508 -22287
rect 8920 -22320 9508 -22304
rect 9938 -22304 9954 -22287
rect 10510 -22287 10712 -22270
rect 10770 -22270 11730 -22232
rect 10770 -22287 10972 -22270
rect 10510 -22304 10526 -22287
rect 9938 -22320 10526 -22304
rect 10956 -22304 10972 -22287
rect 11528 -22287 11730 -22270
rect 11788 -22270 12748 -22232
rect 11788 -22287 11990 -22270
rect 11528 -22304 11544 -22287
rect 10956 -22320 11544 -22304
rect 11974 -22304 11990 -22287
rect 12546 -22287 12748 -22270
rect 12806 -22270 13766 -22232
rect 12806 -22287 13008 -22270
rect 12546 -22304 12562 -22287
rect 11974 -22320 12562 -22304
rect 12992 -22304 13008 -22287
rect 13564 -22287 13766 -22270
rect 13824 -22270 14784 -22232
rect 13824 -22287 14026 -22270
rect 13564 -22304 13580 -22287
rect 12992 -22320 13580 -22304
rect 14010 -22304 14026 -22287
rect 14582 -22287 14784 -22270
rect 14842 -22270 15802 -22232
rect 14842 -22287 15044 -22270
rect 14582 -22304 14598 -22287
rect 14010 -22320 14598 -22304
rect 15028 -22304 15044 -22287
rect 15600 -22287 15802 -22270
rect 15860 -22270 16820 -22232
rect 15860 -22287 16062 -22270
rect 15600 -22304 15616 -22287
rect 15028 -22320 15616 -22304
rect 16046 -22304 16062 -22287
rect 16618 -22287 16820 -22270
rect 16878 -22270 17838 -22232
rect 16878 -22287 17080 -22270
rect 16618 -22304 16634 -22287
rect 16046 -22320 16634 -22304
rect 17064 -22304 17080 -22287
rect 17636 -22287 17838 -22270
rect 17896 -22270 18856 -22232
rect 17896 -22287 18098 -22270
rect 17636 -22304 17652 -22287
rect 17064 -22320 17652 -22304
rect 18082 -22304 18098 -22287
rect 18654 -22287 18856 -22270
rect 18914 -22270 19874 -22232
rect 18914 -22287 19116 -22270
rect 18654 -22304 18670 -22287
rect 18082 -22320 18670 -22304
rect 19100 -22304 19116 -22287
rect 19672 -22287 19874 -22270
rect 19932 -22270 20892 -22232
rect 19932 -22287 20134 -22270
rect 19672 -22304 19688 -22287
rect 19100 -22320 19688 -22304
rect 20118 -22304 20134 -22287
rect 20690 -22287 20892 -22270
rect 20950 -22270 21910 -22232
rect 20950 -22287 21152 -22270
rect 20690 -22304 20706 -22287
rect 20118 -22320 20706 -22304
rect 21136 -22304 21152 -22287
rect 21708 -22287 21910 -22270
rect 21968 -22270 22928 -22232
rect 21968 -22287 22170 -22270
rect 21708 -22304 21724 -22287
rect 21136 -22320 21724 -22304
rect 22154 -22304 22170 -22287
rect 22726 -22287 22928 -22270
rect 22726 -22304 22742 -22287
rect 22154 -22320 22742 -22304
rect 2812 -22792 3400 -22776
rect 2812 -22809 2828 -22792
rect 2626 -22826 2828 -22809
rect 3384 -22809 3400 -22792
rect 3830 -22792 4418 -22776
rect 3830 -22809 3846 -22792
rect 3384 -22826 3586 -22809
rect 2626 -22864 3586 -22826
rect 3644 -22826 3846 -22809
rect 4402 -22809 4418 -22792
rect 4848 -22792 5436 -22776
rect 4848 -22809 4864 -22792
rect 4402 -22826 4604 -22809
rect 3644 -22864 4604 -22826
rect 4662 -22826 4864 -22809
rect 5420 -22809 5436 -22792
rect 5866 -22792 6454 -22776
rect 5866 -22809 5882 -22792
rect 5420 -22826 5622 -22809
rect 4662 -22864 5622 -22826
rect 5680 -22826 5882 -22809
rect 6438 -22809 6454 -22792
rect 6884 -22792 7472 -22776
rect 6884 -22809 6900 -22792
rect 6438 -22826 6640 -22809
rect 5680 -22864 6640 -22826
rect 6698 -22826 6900 -22809
rect 7456 -22809 7472 -22792
rect 7902 -22792 8490 -22776
rect 7902 -22809 7918 -22792
rect 7456 -22826 7658 -22809
rect 6698 -22864 7658 -22826
rect 7716 -22826 7918 -22809
rect 8474 -22809 8490 -22792
rect 8920 -22792 9508 -22776
rect 8920 -22809 8936 -22792
rect 8474 -22826 8676 -22809
rect 7716 -22864 8676 -22826
rect 8734 -22826 8936 -22809
rect 9492 -22809 9508 -22792
rect 9938 -22792 10526 -22776
rect 9938 -22809 9954 -22792
rect 9492 -22826 9694 -22809
rect 8734 -22864 9694 -22826
rect 9752 -22826 9954 -22809
rect 10510 -22809 10526 -22792
rect 10956 -22792 11544 -22776
rect 10956 -22809 10972 -22792
rect 10510 -22826 10712 -22809
rect 9752 -22864 10712 -22826
rect 10770 -22826 10972 -22809
rect 11528 -22809 11544 -22792
rect 11974 -22792 12562 -22776
rect 11974 -22809 11990 -22792
rect 11528 -22826 11730 -22809
rect 10770 -22864 11730 -22826
rect 11788 -22826 11990 -22809
rect 12546 -22809 12562 -22792
rect 12992 -22792 13580 -22776
rect 12992 -22809 13008 -22792
rect 12546 -22826 12748 -22809
rect 11788 -22864 12748 -22826
rect 12806 -22826 13008 -22809
rect 13564 -22809 13580 -22792
rect 14010 -22792 14598 -22776
rect 14010 -22809 14026 -22792
rect 13564 -22826 13766 -22809
rect 12806 -22864 13766 -22826
rect 13824 -22826 14026 -22809
rect 14582 -22809 14598 -22792
rect 15028 -22792 15616 -22776
rect 15028 -22809 15044 -22792
rect 14582 -22826 14784 -22809
rect 13824 -22864 14784 -22826
rect 14842 -22826 15044 -22809
rect 15600 -22809 15616 -22792
rect 16046 -22792 16634 -22776
rect 16046 -22809 16062 -22792
rect 15600 -22826 15802 -22809
rect 14842 -22864 15802 -22826
rect 15860 -22826 16062 -22809
rect 16618 -22809 16634 -22792
rect 17064 -22792 17652 -22776
rect 17064 -22809 17080 -22792
rect 16618 -22826 16820 -22809
rect 15860 -22864 16820 -22826
rect 16878 -22826 17080 -22809
rect 17636 -22809 17652 -22792
rect 18082 -22792 18670 -22776
rect 18082 -22809 18098 -22792
rect 17636 -22826 17838 -22809
rect 16878 -22864 17838 -22826
rect 17896 -22826 18098 -22809
rect 18654 -22809 18670 -22792
rect 19100 -22792 19688 -22776
rect 19100 -22809 19116 -22792
rect 18654 -22826 18856 -22809
rect 17896 -22864 18856 -22826
rect 18914 -22826 19116 -22809
rect 19672 -22809 19688 -22792
rect 20118 -22792 20706 -22776
rect 20118 -22809 20134 -22792
rect 19672 -22826 19874 -22809
rect 18914 -22864 19874 -22826
rect 19932 -22826 20134 -22809
rect 20690 -22809 20706 -22792
rect 21136 -22792 21724 -22776
rect 21136 -22809 21152 -22792
rect 20690 -22826 20892 -22809
rect 19932 -22864 20892 -22826
rect 20950 -22826 21152 -22809
rect 21708 -22809 21724 -22792
rect 22154 -22792 22742 -22776
rect 22154 -22809 22170 -22792
rect 21708 -22826 21910 -22809
rect 20950 -22864 21910 -22826
rect 21968 -22826 22170 -22809
rect 22726 -22809 22742 -22792
rect 22726 -22826 22928 -22809
rect 21968 -22864 22928 -22826
rect 2626 -23502 3586 -23464
rect 2626 -23519 2828 -23502
rect 2812 -23536 2828 -23519
rect 3384 -23519 3586 -23502
rect 3644 -23502 4604 -23464
rect 3644 -23519 3846 -23502
rect 3384 -23536 3400 -23519
rect 2812 -23552 3400 -23536
rect 3830 -23536 3846 -23519
rect 4402 -23519 4604 -23502
rect 4662 -23502 5622 -23464
rect 4662 -23519 4864 -23502
rect 4402 -23536 4418 -23519
rect 3830 -23552 4418 -23536
rect 4848 -23536 4864 -23519
rect 5420 -23519 5622 -23502
rect 5680 -23502 6640 -23464
rect 5680 -23519 5882 -23502
rect 5420 -23536 5436 -23519
rect 4848 -23552 5436 -23536
rect 5866 -23536 5882 -23519
rect 6438 -23519 6640 -23502
rect 6698 -23502 7658 -23464
rect 6698 -23519 6900 -23502
rect 6438 -23536 6454 -23519
rect 5866 -23552 6454 -23536
rect 6884 -23536 6900 -23519
rect 7456 -23519 7658 -23502
rect 7716 -23502 8676 -23464
rect 7716 -23519 7918 -23502
rect 7456 -23536 7472 -23519
rect 6884 -23552 7472 -23536
rect 7902 -23536 7918 -23519
rect 8474 -23519 8676 -23502
rect 8734 -23502 9694 -23464
rect 8734 -23519 8936 -23502
rect 8474 -23536 8490 -23519
rect 7902 -23552 8490 -23536
rect 8920 -23536 8936 -23519
rect 9492 -23519 9694 -23502
rect 9752 -23502 10712 -23464
rect 9752 -23519 9954 -23502
rect 9492 -23536 9508 -23519
rect 8920 -23552 9508 -23536
rect 9938 -23536 9954 -23519
rect 10510 -23519 10712 -23502
rect 10770 -23502 11730 -23464
rect 10770 -23519 10972 -23502
rect 10510 -23536 10526 -23519
rect 9938 -23552 10526 -23536
rect 10956 -23536 10972 -23519
rect 11528 -23519 11730 -23502
rect 11788 -23502 12748 -23464
rect 11788 -23519 11990 -23502
rect 11528 -23536 11544 -23519
rect 10956 -23552 11544 -23536
rect 11974 -23536 11990 -23519
rect 12546 -23519 12748 -23502
rect 12806 -23502 13766 -23464
rect 12806 -23519 13008 -23502
rect 12546 -23536 12562 -23519
rect 11974 -23552 12562 -23536
rect 12992 -23536 13008 -23519
rect 13564 -23519 13766 -23502
rect 13824 -23502 14784 -23464
rect 13824 -23519 14026 -23502
rect 13564 -23536 13580 -23519
rect 12992 -23552 13580 -23536
rect 14010 -23536 14026 -23519
rect 14582 -23519 14784 -23502
rect 14842 -23502 15802 -23464
rect 14842 -23519 15044 -23502
rect 14582 -23536 14598 -23519
rect 14010 -23552 14598 -23536
rect 15028 -23536 15044 -23519
rect 15600 -23519 15802 -23502
rect 15860 -23502 16820 -23464
rect 15860 -23519 16062 -23502
rect 15600 -23536 15616 -23519
rect 15028 -23552 15616 -23536
rect 16046 -23536 16062 -23519
rect 16618 -23519 16820 -23502
rect 16878 -23502 17838 -23464
rect 16878 -23519 17080 -23502
rect 16618 -23536 16634 -23519
rect 16046 -23552 16634 -23536
rect 17064 -23536 17080 -23519
rect 17636 -23519 17838 -23502
rect 17896 -23502 18856 -23464
rect 17896 -23519 18098 -23502
rect 17636 -23536 17652 -23519
rect 17064 -23552 17652 -23536
rect 18082 -23536 18098 -23519
rect 18654 -23519 18856 -23502
rect 18914 -23502 19874 -23464
rect 18914 -23519 19116 -23502
rect 18654 -23536 18670 -23519
rect 18082 -23552 18670 -23536
rect 19100 -23536 19116 -23519
rect 19672 -23519 19874 -23502
rect 19932 -23502 20892 -23464
rect 19932 -23519 20134 -23502
rect 19672 -23536 19688 -23519
rect 19100 -23552 19688 -23536
rect 20118 -23536 20134 -23519
rect 20690 -23519 20892 -23502
rect 20950 -23502 21910 -23464
rect 20950 -23519 21152 -23502
rect 20690 -23536 20706 -23519
rect 20118 -23552 20706 -23536
rect 21136 -23536 21152 -23519
rect 21708 -23519 21910 -23502
rect 21968 -23502 22928 -23464
rect 21968 -23519 22170 -23502
rect 21708 -23536 21724 -23519
rect 21136 -23552 21724 -23536
rect 22154 -23536 22170 -23519
rect 22726 -23519 22928 -23502
rect 22726 -23536 22742 -23519
rect 22154 -23552 22742 -23536
rect 2812 -24026 3400 -24010
rect 2812 -24043 2828 -24026
rect 2626 -24060 2828 -24043
rect 3384 -24043 3400 -24026
rect 3830 -24026 4418 -24010
rect 3830 -24043 3846 -24026
rect 3384 -24060 3586 -24043
rect 2626 -24098 3586 -24060
rect 3644 -24060 3846 -24043
rect 4402 -24043 4418 -24026
rect 4848 -24026 5436 -24010
rect 4848 -24043 4864 -24026
rect 4402 -24060 4604 -24043
rect 3644 -24098 4604 -24060
rect 4662 -24060 4864 -24043
rect 5420 -24043 5436 -24026
rect 5866 -24026 6454 -24010
rect 5866 -24043 5882 -24026
rect 5420 -24060 5622 -24043
rect 4662 -24098 5622 -24060
rect 5680 -24060 5882 -24043
rect 6438 -24043 6454 -24026
rect 6884 -24026 7472 -24010
rect 6884 -24043 6900 -24026
rect 6438 -24060 6640 -24043
rect 5680 -24098 6640 -24060
rect 6698 -24060 6900 -24043
rect 7456 -24043 7472 -24026
rect 7902 -24026 8490 -24010
rect 7902 -24043 7918 -24026
rect 7456 -24060 7658 -24043
rect 6698 -24098 7658 -24060
rect 7716 -24060 7918 -24043
rect 8474 -24043 8490 -24026
rect 8920 -24026 9508 -24010
rect 8920 -24043 8936 -24026
rect 8474 -24060 8676 -24043
rect 7716 -24098 8676 -24060
rect 8734 -24060 8936 -24043
rect 9492 -24043 9508 -24026
rect 9938 -24026 10526 -24010
rect 9938 -24043 9954 -24026
rect 9492 -24060 9694 -24043
rect 8734 -24098 9694 -24060
rect 9752 -24060 9954 -24043
rect 10510 -24043 10526 -24026
rect 10956 -24026 11544 -24010
rect 10956 -24043 10972 -24026
rect 10510 -24060 10712 -24043
rect 9752 -24098 10712 -24060
rect 10770 -24060 10972 -24043
rect 11528 -24043 11544 -24026
rect 11974 -24026 12562 -24010
rect 11974 -24043 11990 -24026
rect 11528 -24060 11730 -24043
rect 10770 -24098 11730 -24060
rect 11788 -24060 11990 -24043
rect 12546 -24043 12562 -24026
rect 12992 -24026 13580 -24010
rect 12992 -24043 13008 -24026
rect 12546 -24060 12748 -24043
rect 11788 -24098 12748 -24060
rect 12806 -24060 13008 -24043
rect 13564 -24043 13580 -24026
rect 14010 -24026 14598 -24010
rect 14010 -24043 14026 -24026
rect 13564 -24060 13766 -24043
rect 12806 -24098 13766 -24060
rect 13824 -24060 14026 -24043
rect 14582 -24043 14598 -24026
rect 15028 -24026 15616 -24010
rect 15028 -24043 15044 -24026
rect 14582 -24060 14784 -24043
rect 13824 -24098 14784 -24060
rect 14842 -24060 15044 -24043
rect 15600 -24043 15616 -24026
rect 16046 -24026 16634 -24010
rect 16046 -24043 16062 -24026
rect 15600 -24060 15802 -24043
rect 14842 -24098 15802 -24060
rect 15860 -24060 16062 -24043
rect 16618 -24043 16634 -24026
rect 17064 -24026 17652 -24010
rect 17064 -24043 17080 -24026
rect 16618 -24060 16820 -24043
rect 15860 -24098 16820 -24060
rect 16878 -24060 17080 -24043
rect 17636 -24043 17652 -24026
rect 18082 -24026 18670 -24010
rect 18082 -24043 18098 -24026
rect 17636 -24060 17838 -24043
rect 16878 -24098 17838 -24060
rect 17896 -24060 18098 -24043
rect 18654 -24043 18670 -24026
rect 19100 -24026 19688 -24010
rect 19100 -24043 19116 -24026
rect 18654 -24060 18856 -24043
rect 17896 -24098 18856 -24060
rect 18914 -24060 19116 -24043
rect 19672 -24043 19688 -24026
rect 20118 -24026 20706 -24010
rect 20118 -24043 20134 -24026
rect 19672 -24060 19874 -24043
rect 18914 -24098 19874 -24060
rect 19932 -24060 20134 -24043
rect 20690 -24043 20706 -24026
rect 21136 -24026 21724 -24010
rect 21136 -24043 21152 -24026
rect 20690 -24060 20892 -24043
rect 19932 -24098 20892 -24060
rect 20950 -24060 21152 -24043
rect 21708 -24043 21724 -24026
rect 22154 -24026 22742 -24010
rect 22154 -24043 22170 -24026
rect 21708 -24060 21910 -24043
rect 20950 -24098 21910 -24060
rect 21968 -24060 22170 -24043
rect 22726 -24043 22742 -24026
rect 22726 -24060 22928 -24043
rect 21968 -24098 22928 -24060
rect 2626 -24736 3586 -24698
rect 2626 -24753 2828 -24736
rect 2812 -24770 2828 -24753
rect 3384 -24753 3586 -24736
rect 3644 -24736 4604 -24698
rect 3644 -24753 3846 -24736
rect 3384 -24770 3400 -24753
rect 2812 -24786 3400 -24770
rect 3830 -24770 3846 -24753
rect 4402 -24753 4604 -24736
rect 4662 -24736 5622 -24698
rect 4662 -24753 4864 -24736
rect 4402 -24770 4418 -24753
rect 3830 -24786 4418 -24770
rect 4848 -24770 4864 -24753
rect 5420 -24753 5622 -24736
rect 5680 -24736 6640 -24698
rect 5680 -24753 5882 -24736
rect 5420 -24770 5436 -24753
rect 4848 -24786 5436 -24770
rect 5866 -24770 5882 -24753
rect 6438 -24753 6640 -24736
rect 6698 -24736 7658 -24698
rect 6698 -24753 6900 -24736
rect 6438 -24770 6454 -24753
rect 5866 -24786 6454 -24770
rect 6884 -24770 6900 -24753
rect 7456 -24753 7658 -24736
rect 7716 -24736 8676 -24698
rect 7716 -24753 7918 -24736
rect 7456 -24770 7472 -24753
rect 6884 -24786 7472 -24770
rect 7902 -24770 7918 -24753
rect 8474 -24753 8676 -24736
rect 8734 -24736 9694 -24698
rect 8734 -24753 8936 -24736
rect 8474 -24770 8490 -24753
rect 7902 -24786 8490 -24770
rect 8920 -24770 8936 -24753
rect 9492 -24753 9694 -24736
rect 9752 -24736 10712 -24698
rect 9752 -24753 9954 -24736
rect 9492 -24770 9508 -24753
rect 8920 -24786 9508 -24770
rect 9938 -24770 9954 -24753
rect 10510 -24753 10712 -24736
rect 10770 -24736 11730 -24698
rect 10770 -24753 10972 -24736
rect 10510 -24770 10526 -24753
rect 9938 -24786 10526 -24770
rect 10956 -24770 10972 -24753
rect 11528 -24753 11730 -24736
rect 11788 -24736 12748 -24698
rect 11788 -24753 11990 -24736
rect 11528 -24770 11544 -24753
rect 10956 -24786 11544 -24770
rect 11974 -24770 11990 -24753
rect 12546 -24753 12748 -24736
rect 12806 -24736 13766 -24698
rect 12806 -24753 13008 -24736
rect 12546 -24770 12562 -24753
rect 11974 -24786 12562 -24770
rect 12992 -24770 13008 -24753
rect 13564 -24753 13766 -24736
rect 13824 -24736 14784 -24698
rect 13824 -24753 14026 -24736
rect 13564 -24770 13580 -24753
rect 12992 -24786 13580 -24770
rect 14010 -24770 14026 -24753
rect 14582 -24753 14784 -24736
rect 14842 -24736 15802 -24698
rect 14842 -24753 15044 -24736
rect 14582 -24770 14598 -24753
rect 14010 -24786 14598 -24770
rect 15028 -24770 15044 -24753
rect 15600 -24753 15802 -24736
rect 15860 -24736 16820 -24698
rect 15860 -24753 16062 -24736
rect 15600 -24770 15616 -24753
rect 15028 -24786 15616 -24770
rect 16046 -24770 16062 -24753
rect 16618 -24753 16820 -24736
rect 16878 -24736 17838 -24698
rect 16878 -24753 17080 -24736
rect 16618 -24770 16634 -24753
rect 16046 -24786 16634 -24770
rect 17064 -24770 17080 -24753
rect 17636 -24753 17838 -24736
rect 17896 -24736 18856 -24698
rect 17896 -24753 18098 -24736
rect 17636 -24770 17652 -24753
rect 17064 -24786 17652 -24770
rect 18082 -24770 18098 -24753
rect 18654 -24753 18856 -24736
rect 18914 -24736 19874 -24698
rect 18914 -24753 19116 -24736
rect 18654 -24770 18670 -24753
rect 18082 -24786 18670 -24770
rect 19100 -24770 19116 -24753
rect 19672 -24753 19874 -24736
rect 19932 -24736 20892 -24698
rect 19932 -24753 20134 -24736
rect 19672 -24770 19688 -24753
rect 19100 -24786 19688 -24770
rect 20118 -24770 20134 -24753
rect 20690 -24753 20892 -24736
rect 20950 -24736 21910 -24698
rect 20950 -24753 21152 -24736
rect 20690 -24770 20706 -24753
rect 20118 -24786 20706 -24770
rect 21136 -24770 21152 -24753
rect 21708 -24753 21910 -24736
rect 21968 -24736 22928 -24698
rect 21968 -24753 22170 -24736
rect 21708 -24770 21724 -24753
rect 21136 -24786 21724 -24770
rect 22154 -24770 22170 -24753
rect 22726 -24753 22928 -24736
rect 22726 -24770 22742 -24753
rect 22154 -24786 22742 -24770
<< polycont >>
rect -8936 -12474 -8380 -12440
rect -7918 -12474 -7362 -12440
rect -6900 -12474 -6344 -12440
rect -5882 -12474 -5326 -12440
rect -4864 -12474 -4308 -12440
rect -3846 -12474 -3290 -12440
rect -2828 -12474 -2272 -12440
rect -1810 -12474 -1254 -12440
rect -792 -12474 -236 -12440
rect -8936 -13184 -8380 -13150
rect -7918 -13184 -7362 -13150
rect -6900 -13184 -6344 -13150
rect -5882 -13184 -5326 -13150
rect -4864 -13184 -4308 -13150
rect -3846 -13184 -3290 -13150
rect -2828 -13184 -2272 -13150
rect -1810 -13184 -1254 -13150
rect -792 -13184 -236 -13150
rect -8936 -13292 -8380 -13258
rect -7918 -13292 -7362 -13258
rect -6900 -13292 -6344 -13258
rect -5882 -13292 -5326 -13258
rect -4864 -13292 -4308 -13258
rect -3846 -13292 -3290 -13258
rect -2828 -13292 -2272 -13258
rect -1810 -13292 -1254 -13258
rect -792 -13292 -236 -13258
rect -8936 -14002 -8380 -13968
rect -7918 -14002 -7362 -13968
rect -6900 -14002 -6344 -13968
rect -5882 -14002 -5326 -13968
rect -4864 -14002 -4308 -13968
rect -3846 -14002 -3290 -13968
rect -2828 -14002 -2272 -13968
rect -1810 -14002 -1254 -13968
rect -792 -14002 -236 -13968
rect -8936 -14110 -8380 -14076
rect -7918 -14110 -7362 -14076
rect -6900 -14110 -6344 -14076
rect -5882 -14110 -5326 -14076
rect -4864 -14110 -4308 -14076
rect -3846 -14110 -3290 -14076
rect -2828 -14110 -2272 -14076
rect -1810 -14110 -1254 -14076
rect -792 -14110 -236 -14076
rect 2830 -14194 3386 -14160
rect 3848 -14194 4404 -14160
rect 4866 -14194 5422 -14160
rect 5884 -14194 6440 -14160
rect 6902 -14194 7458 -14160
rect 7920 -14194 8476 -14160
rect 8938 -14194 9494 -14160
rect 9956 -14194 10512 -14160
rect 10974 -14194 11530 -14160
rect 11992 -14194 12548 -14160
rect 13010 -14194 13566 -14160
rect 14028 -14194 14584 -14160
rect 15046 -14194 15602 -14160
rect 16064 -14194 16620 -14160
rect 17082 -14194 17638 -14160
rect 18100 -14194 18656 -14160
rect 19118 -14194 19674 -14160
rect 20136 -14194 20692 -14160
rect 21154 -14194 21710 -14160
rect 22172 -14194 22728 -14160
rect -8936 -14820 -8380 -14786
rect -7918 -14820 -7362 -14786
rect -6900 -14820 -6344 -14786
rect -5882 -14820 -5326 -14786
rect -4864 -14820 -4308 -14786
rect -3846 -14820 -3290 -14786
rect -2828 -14820 -2272 -14786
rect -1810 -14820 -1254 -14786
rect -792 -14820 -236 -14786
rect -8936 -14928 -8380 -14894
rect -7918 -14928 -7362 -14894
rect -6900 -14928 -6344 -14894
rect -5882 -14928 -5326 -14894
rect -4864 -14928 -4308 -14894
rect -3846 -14928 -3290 -14894
rect -2828 -14928 -2272 -14894
rect -1810 -14928 -1254 -14894
rect -792 -14928 -236 -14894
rect 2830 -14904 3386 -14870
rect 3848 -14904 4404 -14870
rect 4866 -14904 5422 -14870
rect 5884 -14904 6440 -14870
rect 6902 -14904 7458 -14870
rect 7920 -14904 8476 -14870
rect 8938 -14904 9494 -14870
rect 9956 -14904 10512 -14870
rect 10974 -14904 11530 -14870
rect 11992 -14904 12548 -14870
rect 13010 -14904 13566 -14870
rect 14028 -14904 14584 -14870
rect 15046 -14904 15602 -14870
rect 16064 -14904 16620 -14870
rect 17082 -14904 17638 -14870
rect 18100 -14904 18656 -14870
rect 19118 -14904 19674 -14870
rect 20136 -14904 20692 -14870
rect 21154 -14904 21710 -14870
rect 22172 -14904 22728 -14870
rect 2830 -15426 3386 -15392
rect 3848 -15426 4404 -15392
rect 4866 -15426 5422 -15392
rect 5884 -15426 6440 -15392
rect 6902 -15426 7458 -15392
rect 7920 -15426 8476 -15392
rect 8938 -15426 9494 -15392
rect 9956 -15426 10512 -15392
rect 10974 -15426 11530 -15392
rect 11992 -15426 12548 -15392
rect 13010 -15426 13566 -15392
rect 14028 -15426 14584 -15392
rect 15046 -15426 15602 -15392
rect 16064 -15426 16620 -15392
rect 17082 -15426 17638 -15392
rect 18100 -15426 18656 -15392
rect 19118 -15426 19674 -15392
rect 20136 -15426 20692 -15392
rect 21154 -15426 21710 -15392
rect 22172 -15426 22728 -15392
rect -8936 -15638 -8380 -15604
rect -7918 -15638 -7362 -15604
rect -6900 -15638 -6344 -15604
rect -5882 -15638 -5326 -15604
rect -4864 -15638 -4308 -15604
rect -3846 -15638 -3290 -15604
rect -2828 -15638 -2272 -15604
rect -1810 -15638 -1254 -15604
rect -792 -15638 -236 -15604
rect -8936 -15746 -8380 -15712
rect -7918 -15746 -7362 -15712
rect -6900 -15746 -6344 -15712
rect -5882 -15746 -5326 -15712
rect -4864 -15746 -4308 -15712
rect -3846 -15746 -3290 -15712
rect -2828 -15746 -2272 -15712
rect -1810 -15746 -1254 -15712
rect -792 -15746 -236 -15712
rect 2830 -16136 3386 -16102
rect 3848 -16136 4404 -16102
rect 4866 -16136 5422 -16102
rect 5884 -16136 6440 -16102
rect 6902 -16136 7458 -16102
rect 7920 -16136 8476 -16102
rect 8938 -16136 9494 -16102
rect 9956 -16136 10512 -16102
rect 10974 -16136 11530 -16102
rect 11992 -16136 12548 -16102
rect 13010 -16136 13566 -16102
rect 14028 -16136 14584 -16102
rect 15046 -16136 15602 -16102
rect 16064 -16136 16620 -16102
rect 17082 -16136 17638 -16102
rect 18100 -16136 18656 -16102
rect 19118 -16136 19674 -16102
rect 20136 -16136 20692 -16102
rect 21154 -16136 21710 -16102
rect 22172 -16136 22728 -16102
rect -8936 -16456 -8380 -16422
rect -7918 -16456 -7362 -16422
rect -6900 -16456 -6344 -16422
rect -5882 -16456 -5326 -16422
rect -4864 -16456 -4308 -16422
rect -3846 -16456 -3290 -16422
rect -2828 -16456 -2272 -16422
rect -1810 -16456 -1254 -16422
rect -792 -16456 -236 -16422
rect -8936 -16564 -8380 -16530
rect -7918 -16564 -7362 -16530
rect -6900 -16564 -6344 -16530
rect -5882 -16564 -5326 -16530
rect -4864 -16564 -4308 -16530
rect -3846 -16564 -3290 -16530
rect -2828 -16564 -2272 -16530
rect -1810 -16564 -1254 -16530
rect -792 -16564 -236 -16530
rect 2828 -16660 3384 -16626
rect 3846 -16660 4402 -16626
rect 4864 -16660 5420 -16626
rect 5882 -16660 6438 -16626
rect 6900 -16660 7456 -16626
rect 7918 -16660 8474 -16626
rect 8936 -16660 9492 -16626
rect 9954 -16660 10510 -16626
rect 10972 -16660 11528 -16626
rect 11990 -16660 12546 -16626
rect 13008 -16660 13564 -16626
rect 14026 -16660 14582 -16626
rect 15044 -16660 15600 -16626
rect 16062 -16660 16618 -16626
rect 17080 -16660 17636 -16626
rect 18098 -16660 18654 -16626
rect 19116 -16660 19672 -16626
rect 20134 -16660 20690 -16626
rect 21152 -16660 21708 -16626
rect 22170 -16660 22726 -16626
rect -8936 -17274 -8380 -17240
rect -7918 -17274 -7362 -17240
rect -6900 -17274 -6344 -17240
rect -5882 -17274 -5326 -17240
rect -4864 -17274 -4308 -17240
rect -3846 -17274 -3290 -17240
rect -2828 -17274 -2272 -17240
rect -1810 -17274 -1254 -17240
rect -792 -17274 -236 -17240
rect -8936 -17382 -8380 -17348
rect -7918 -17382 -7362 -17348
rect -6900 -17382 -6344 -17348
rect -5882 -17382 -5326 -17348
rect -4864 -17382 -4308 -17348
rect -3846 -17382 -3290 -17348
rect -2828 -17382 -2272 -17348
rect -1810 -17382 -1254 -17348
rect -792 -17382 -236 -17348
rect 2828 -17370 3384 -17336
rect 3846 -17370 4402 -17336
rect 4864 -17370 5420 -17336
rect 5882 -17370 6438 -17336
rect 6900 -17370 7456 -17336
rect 7918 -17370 8474 -17336
rect 8936 -17370 9492 -17336
rect 9954 -17370 10510 -17336
rect 10972 -17370 11528 -17336
rect 11990 -17370 12546 -17336
rect 13008 -17370 13564 -17336
rect 14026 -17370 14582 -17336
rect 15044 -17370 15600 -17336
rect 16062 -17370 16618 -17336
rect 17080 -17370 17636 -17336
rect 18098 -17370 18654 -17336
rect 19116 -17370 19672 -17336
rect 20134 -17370 20690 -17336
rect 21152 -17370 21708 -17336
rect 22170 -17370 22726 -17336
rect 2828 -17894 3384 -17860
rect 3846 -17894 4402 -17860
rect 4864 -17894 5420 -17860
rect 5882 -17894 6438 -17860
rect 6900 -17894 7456 -17860
rect 7918 -17894 8474 -17860
rect 8936 -17894 9492 -17860
rect 9954 -17894 10510 -17860
rect 10972 -17894 11528 -17860
rect 11990 -17894 12546 -17860
rect 13008 -17894 13564 -17860
rect 14026 -17894 14582 -17860
rect 15044 -17894 15600 -17860
rect 16062 -17894 16618 -17860
rect 17080 -17894 17636 -17860
rect 18098 -17894 18654 -17860
rect 19116 -17894 19672 -17860
rect 20134 -17894 20690 -17860
rect 21152 -17894 21708 -17860
rect 22170 -17894 22726 -17860
rect -8936 -18092 -8380 -18058
rect -7918 -18092 -7362 -18058
rect -6900 -18092 -6344 -18058
rect -5882 -18092 -5326 -18058
rect -4864 -18092 -4308 -18058
rect -3846 -18092 -3290 -18058
rect -2828 -18092 -2272 -18058
rect -1810 -18092 -1254 -18058
rect -792 -18092 -236 -18058
rect -8936 -18200 -8380 -18166
rect -7918 -18200 -7362 -18166
rect -6900 -18200 -6344 -18166
rect -5882 -18200 -5326 -18166
rect -4864 -18200 -4308 -18166
rect -3846 -18200 -3290 -18166
rect -2828 -18200 -2272 -18166
rect -1810 -18200 -1254 -18166
rect -792 -18200 -236 -18166
rect 2828 -18604 3384 -18570
rect 3846 -18604 4402 -18570
rect 4864 -18604 5420 -18570
rect 5882 -18604 6438 -18570
rect 6900 -18604 7456 -18570
rect 7918 -18604 8474 -18570
rect 8936 -18604 9492 -18570
rect 9954 -18604 10510 -18570
rect 10972 -18604 11528 -18570
rect 11990 -18604 12546 -18570
rect 13008 -18604 13564 -18570
rect 14026 -18604 14582 -18570
rect 15044 -18604 15600 -18570
rect 16062 -18604 16618 -18570
rect 17080 -18604 17636 -18570
rect 18098 -18604 18654 -18570
rect 19116 -18604 19672 -18570
rect 20134 -18604 20690 -18570
rect 21152 -18604 21708 -18570
rect 22170 -18604 22726 -18570
rect -8936 -18910 -8380 -18876
rect -7918 -18910 -7362 -18876
rect -6900 -18910 -6344 -18876
rect -5882 -18910 -5326 -18876
rect -4864 -18910 -4308 -18876
rect -3846 -18910 -3290 -18876
rect -2828 -18910 -2272 -18876
rect -1810 -18910 -1254 -18876
rect -792 -18910 -236 -18876
rect 2828 -19126 3384 -19092
rect 3846 -19126 4402 -19092
rect 4864 -19126 5420 -19092
rect 5882 -19126 6438 -19092
rect 6900 -19126 7456 -19092
rect 7918 -19126 8474 -19092
rect 8936 -19126 9492 -19092
rect 9954 -19126 10510 -19092
rect 10972 -19126 11528 -19092
rect 11990 -19126 12546 -19092
rect 13008 -19126 13564 -19092
rect 14026 -19126 14582 -19092
rect 15044 -19126 15600 -19092
rect 16062 -19126 16618 -19092
rect 17080 -19126 17636 -19092
rect 18098 -19126 18654 -19092
rect 19116 -19126 19672 -19092
rect 20134 -19126 20690 -19092
rect 21152 -19126 21708 -19092
rect 22170 -19126 22726 -19092
rect 2828 -19836 3384 -19802
rect 3846 -19836 4402 -19802
rect 4864 -19836 5420 -19802
rect 5882 -19836 6438 -19802
rect 6900 -19836 7456 -19802
rect 7918 -19836 8474 -19802
rect 8936 -19836 9492 -19802
rect 9954 -19836 10510 -19802
rect 10972 -19836 11528 -19802
rect 11990 -19836 12546 -19802
rect 13008 -19836 13564 -19802
rect 14026 -19836 14582 -19802
rect 15044 -19836 15600 -19802
rect 16062 -19836 16618 -19802
rect 17080 -19836 17636 -19802
rect 18098 -19836 18654 -19802
rect 19116 -19836 19672 -19802
rect 20134 -19836 20690 -19802
rect 21152 -19836 21708 -19802
rect 22170 -19836 22726 -19802
rect 2828 -20360 3384 -20326
rect 3846 -20360 4402 -20326
rect 4864 -20360 5420 -20326
rect 5882 -20360 6438 -20326
rect 6900 -20360 7456 -20326
rect 7918 -20360 8474 -20326
rect 8936 -20360 9492 -20326
rect 9954 -20360 10510 -20326
rect 10972 -20360 11528 -20326
rect 11990 -20360 12546 -20326
rect 13008 -20360 13564 -20326
rect 14026 -20360 14582 -20326
rect 15044 -20360 15600 -20326
rect 16062 -20360 16618 -20326
rect 17080 -20360 17636 -20326
rect 18098 -20360 18654 -20326
rect 19116 -20360 19672 -20326
rect 20134 -20360 20690 -20326
rect 21152 -20360 21708 -20326
rect 22170 -20360 22726 -20326
rect 2828 -21070 3384 -21036
rect 3846 -21070 4402 -21036
rect 4864 -21070 5420 -21036
rect 5882 -21070 6438 -21036
rect 6900 -21070 7456 -21036
rect 7918 -21070 8474 -21036
rect 8936 -21070 9492 -21036
rect 9954 -21070 10510 -21036
rect 10972 -21070 11528 -21036
rect 11990 -21070 12546 -21036
rect 13008 -21070 13564 -21036
rect 14026 -21070 14582 -21036
rect 15044 -21070 15600 -21036
rect 16062 -21070 16618 -21036
rect 17080 -21070 17636 -21036
rect 18098 -21070 18654 -21036
rect 19116 -21070 19672 -21036
rect 20134 -21070 20690 -21036
rect 21152 -21070 21708 -21036
rect 22170 -21070 22726 -21036
rect 2828 -21594 3384 -21560
rect 3846 -21594 4402 -21560
rect 4864 -21594 5420 -21560
rect 5882 -21594 6438 -21560
rect 6900 -21594 7456 -21560
rect 7918 -21594 8474 -21560
rect 8936 -21594 9492 -21560
rect 9954 -21594 10510 -21560
rect 10972 -21594 11528 -21560
rect 11990 -21594 12546 -21560
rect 13008 -21594 13564 -21560
rect 14026 -21594 14582 -21560
rect 15044 -21594 15600 -21560
rect 16062 -21594 16618 -21560
rect 17080 -21594 17636 -21560
rect 18098 -21594 18654 -21560
rect 19116 -21594 19672 -21560
rect 20134 -21594 20690 -21560
rect 21152 -21594 21708 -21560
rect 22170 -21594 22726 -21560
rect 2828 -22304 3384 -22270
rect 3846 -22304 4402 -22270
rect 4864 -22304 5420 -22270
rect 5882 -22304 6438 -22270
rect 6900 -22304 7456 -22270
rect 7918 -22304 8474 -22270
rect 8936 -22304 9492 -22270
rect 9954 -22304 10510 -22270
rect 10972 -22304 11528 -22270
rect 11990 -22304 12546 -22270
rect 13008 -22304 13564 -22270
rect 14026 -22304 14582 -22270
rect 15044 -22304 15600 -22270
rect 16062 -22304 16618 -22270
rect 17080 -22304 17636 -22270
rect 18098 -22304 18654 -22270
rect 19116 -22304 19672 -22270
rect 20134 -22304 20690 -22270
rect 21152 -22304 21708 -22270
rect 22170 -22304 22726 -22270
rect 2828 -22826 3384 -22792
rect 3846 -22826 4402 -22792
rect 4864 -22826 5420 -22792
rect 5882 -22826 6438 -22792
rect 6900 -22826 7456 -22792
rect 7918 -22826 8474 -22792
rect 8936 -22826 9492 -22792
rect 9954 -22826 10510 -22792
rect 10972 -22826 11528 -22792
rect 11990 -22826 12546 -22792
rect 13008 -22826 13564 -22792
rect 14026 -22826 14582 -22792
rect 15044 -22826 15600 -22792
rect 16062 -22826 16618 -22792
rect 17080 -22826 17636 -22792
rect 18098 -22826 18654 -22792
rect 19116 -22826 19672 -22792
rect 20134 -22826 20690 -22792
rect 21152 -22826 21708 -22792
rect 22170 -22826 22726 -22792
rect 2828 -23536 3384 -23502
rect 3846 -23536 4402 -23502
rect 4864 -23536 5420 -23502
rect 5882 -23536 6438 -23502
rect 6900 -23536 7456 -23502
rect 7918 -23536 8474 -23502
rect 8936 -23536 9492 -23502
rect 9954 -23536 10510 -23502
rect 10972 -23536 11528 -23502
rect 11990 -23536 12546 -23502
rect 13008 -23536 13564 -23502
rect 14026 -23536 14582 -23502
rect 15044 -23536 15600 -23502
rect 16062 -23536 16618 -23502
rect 17080 -23536 17636 -23502
rect 18098 -23536 18654 -23502
rect 19116 -23536 19672 -23502
rect 20134 -23536 20690 -23502
rect 21152 -23536 21708 -23502
rect 22170 -23536 22726 -23502
rect 2828 -24060 3384 -24026
rect 3846 -24060 4402 -24026
rect 4864 -24060 5420 -24026
rect 5882 -24060 6438 -24026
rect 6900 -24060 7456 -24026
rect 7918 -24060 8474 -24026
rect 8936 -24060 9492 -24026
rect 9954 -24060 10510 -24026
rect 10972 -24060 11528 -24026
rect 11990 -24060 12546 -24026
rect 13008 -24060 13564 -24026
rect 14026 -24060 14582 -24026
rect 15044 -24060 15600 -24026
rect 16062 -24060 16618 -24026
rect 17080 -24060 17636 -24026
rect 18098 -24060 18654 -24026
rect 19116 -24060 19672 -24026
rect 20134 -24060 20690 -24026
rect 21152 -24060 21708 -24026
rect 22170 -24060 22726 -24026
rect 2828 -24770 3384 -24736
rect 3846 -24770 4402 -24736
rect 4864 -24770 5420 -24736
rect 5882 -24770 6438 -24736
rect 6900 -24770 7456 -24736
rect 7918 -24770 8474 -24736
rect 8936 -24770 9492 -24736
rect 9954 -24770 10510 -24736
rect 10972 -24770 11528 -24736
rect 11990 -24770 12546 -24736
rect 13008 -24770 13564 -24736
rect 14026 -24770 14582 -24736
rect 15044 -24770 15600 -24736
rect 16062 -24770 16618 -24736
rect 17080 -24770 17636 -24736
rect 18098 -24770 18654 -24736
rect 19116 -24770 19672 -24736
rect 20134 -24770 20690 -24736
rect 21152 -24770 21708 -24736
rect 22170 -24770 22726 -24736
<< locali >>
rect 378 4160 478 4322
rect 378 -10348 478 -10186
rect 24722 4160 24822 4322
rect 24722 -10348 24822 -10186
rect -12322 -11340 -12222 -11178
rect 24822 -11340 24922 -11178
rect -8952 -12474 -8936 -12440
rect -8380 -12474 -8364 -12440
rect -7934 -12474 -7918 -12440
rect -7362 -12474 -7346 -12440
rect -6916 -12474 -6900 -12440
rect -6344 -12474 -6328 -12440
rect -5898 -12474 -5882 -12440
rect -5326 -12474 -5310 -12440
rect -4880 -12474 -4864 -12440
rect -4308 -12474 -4292 -12440
rect -3862 -12474 -3846 -12440
rect -3290 -12474 -3274 -12440
rect -2844 -12474 -2828 -12440
rect -2272 -12474 -2256 -12440
rect -1826 -12474 -1810 -12440
rect -1254 -12474 -1238 -12440
rect -808 -12474 -792 -12440
rect -236 -12474 -220 -12440
rect -9184 -12524 -9150 -12508
rect -9184 -13116 -9150 -13100
rect -8166 -12524 -8132 -12508
rect -8166 -13116 -8132 -13100
rect -7148 -12524 -7114 -12508
rect -7148 -13116 -7114 -13100
rect -6130 -12524 -6096 -12508
rect -6130 -13116 -6096 -13100
rect -5112 -12524 -5078 -12508
rect -5112 -13116 -5078 -13100
rect -4094 -12524 -4060 -12508
rect -4094 -13116 -4060 -13100
rect -3076 -12524 -3042 -12508
rect -3076 -13116 -3042 -13100
rect -2058 -12524 -2024 -12508
rect -2058 -13116 -2024 -13100
rect -1040 -12524 -1006 -12508
rect -1040 -13116 -1006 -13100
rect -22 -12524 12 -12508
rect -22 -13116 12 -13100
rect -8952 -13184 -8936 -13150
rect -8380 -13184 -8364 -13150
rect -7934 -13184 -7918 -13150
rect -7362 -13184 -7346 -13150
rect -6916 -13184 -6900 -13150
rect -6344 -13184 -6328 -13150
rect -5898 -13184 -5882 -13150
rect -5326 -13184 -5310 -13150
rect -4880 -13184 -4864 -13150
rect -4308 -13184 -4292 -13150
rect -3862 -13184 -3846 -13150
rect -3290 -13184 -3274 -13150
rect -2844 -13184 -2828 -13150
rect -2272 -13184 -2256 -13150
rect -1826 -13184 -1810 -13150
rect -1254 -13184 -1238 -13150
rect -808 -13184 -792 -13150
rect -236 -13184 -220 -13150
rect -8952 -13292 -8936 -13258
rect -8380 -13292 -8364 -13258
rect -7934 -13292 -7918 -13258
rect -7362 -13292 -7346 -13258
rect -6916 -13292 -6900 -13258
rect -6344 -13292 -6328 -13258
rect -5898 -13292 -5882 -13258
rect -5326 -13292 -5310 -13258
rect -4880 -13292 -4864 -13258
rect -4308 -13292 -4292 -13258
rect -3862 -13292 -3846 -13258
rect -3290 -13292 -3274 -13258
rect -2844 -13292 -2828 -13258
rect -2272 -13292 -2256 -13258
rect -1826 -13292 -1810 -13258
rect -1254 -13292 -1238 -13258
rect -808 -13292 -792 -13258
rect -236 -13292 -220 -13258
rect -3592 -13294 -3532 -13292
rect -9184 -13342 -9150 -13326
rect -9184 -13934 -9150 -13918
rect -8166 -13342 -8132 -13326
rect -8166 -13934 -8132 -13918
rect -7148 -13342 -7114 -13326
rect -7148 -13934 -7114 -13918
rect -6130 -13342 -6096 -13326
rect -6130 -13934 -6096 -13918
rect -5112 -13342 -5078 -13326
rect -5112 -13934 -5078 -13918
rect -4094 -13342 -4060 -13326
rect -4094 -13934 -4060 -13918
rect -3076 -13342 -3042 -13326
rect -3076 -13934 -3042 -13918
rect -2058 -13342 -2024 -13326
rect -2058 -13934 -2024 -13918
rect -1040 -13342 -1006 -13326
rect -1040 -13934 -1006 -13918
rect -22 -13342 12 -13326
rect -22 -13934 12 -13918
rect -7660 -13968 -7600 -13966
rect -6646 -13968 -6586 -13966
rect -2572 -13968 -2512 -13966
rect -1556 -13968 -1496 -13966
rect -8952 -14002 -8936 -13968
rect -8380 -14002 -8364 -13968
rect -7934 -14002 -7918 -13968
rect -7362 -14002 -7346 -13968
rect -6916 -14002 -6900 -13968
rect -6344 -14002 -6328 -13968
rect -5898 -14002 -5882 -13968
rect -5326 -14002 -5310 -13968
rect -4880 -14002 -4864 -13968
rect -4308 -14002 -4292 -13968
rect -3862 -14002 -3846 -13968
rect -3290 -14002 -3274 -13968
rect -2844 -14002 -2828 -13968
rect -2272 -14002 -2256 -13968
rect -1826 -14002 -1810 -13968
rect -1254 -14002 -1238 -13968
rect -808 -14002 -792 -13968
rect -236 -14002 -220 -13968
rect -8952 -14110 -8936 -14076
rect -8380 -14110 -8364 -14076
rect -7934 -14110 -7918 -14076
rect -7362 -14110 -7346 -14076
rect -6916 -14110 -6900 -14076
rect -6344 -14110 -6328 -14076
rect -5898 -14110 -5882 -14076
rect -5326 -14110 -5310 -14076
rect -4880 -14110 -4864 -14076
rect -4308 -14110 -4292 -14076
rect -3862 -14110 -3846 -14076
rect -3290 -14110 -3274 -14076
rect -2844 -14110 -2828 -14076
rect -2272 -14110 -2256 -14076
rect -1826 -14110 -1810 -14076
rect -1254 -14110 -1238 -14076
rect -808 -14110 -792 -14076
rect -236 -14110 -220 -14076
rect -9184 -14160 -9150 -14144
rect -9184 -14752 -9150 -14736
rect -8166 -14160 -8132 -14144
rect -8166 -14752 -8132 -14736
rect -7148 -14160 -7114 -14144
rect -7148 -14752 -7114 -14736
rect -6130 -14160 -6096 -14144
rect -6130 -14752 -6096 -14736
rect -5112 -14160 -5078 -14144
rect -5112 -14752 -5078 -14736
rect -4094 -14160 -4060 -14144
rect -4094 -14752 -4060 -14736
rect -3076 -14160 -3042 -14144
rect -3076 -14752 -3042 -14736
rect -2058 -14160 -2024 -14144
rect -2058 -14752 -2024 -14736
rect -1040 -14160 -1006 -14144
rect -1040 -14752 -1006 -14736
rect -22 -14160 12 -14144
rect 2814 -14194 2830 -14160
rect 3386 -14194 3402 -14160
rect 3832 -14194 3848 -14160
rect 4404 -14194 4420 -14160
rect 4850 -14194 4866 -14160
rect 5422 -14194 5438 -14160
rect 5868 -14194 5884 -14160
rect 6440 -14194 6456 -14160
rect 6886 -14194 6902 -14160
rect 7458 -14194 7474 -14160
rect 7904 -14194 7920 -14160
rect 8476 -14194 8492 -14160
rect 8922 -14194 8938 -14160
rect 9494 -14194 9510 -14160
rect 9940 -14194 9956 -14160
rect 10512 -14194 10528 -14160
rect 10958 -14194 10974 -14160
rect 11530 -14194 11546 -14160
rect 11976 -14194 11992 -14160
rect 12548 -14194 12564 -14160
rect 12994 -14194 13010 -14160
rect 13566 -14194 13582 -14160
rect 14012 -14194 14028 -14160
rect 14584 -14194 14600 -14160
rect 15030 -14194 15046 -14160
rect 15602 -14194 15618 -14160
rect 16048 -14194 16064 -14160
rect 16620 -14194 16636 -14160
rect 17066 -14194 17082 -14160
rect 17638 -14194 17654 -14160
rect 18084 -14194 18100 -14160
rect 18656 -14194 18672 -14160
rect 19102 -14194 19118 -14160
rect 19674 -14194 19690 -14160
rect 20120 -14194 20136 -14160
rect 20692 -14194 20708 -14160
rect 21138 -14194 21154 -14160
rect 21710 -14194 21726 -14160
rect 22156 -14194 22172 -14160
rect 22728 -14194 22744 -14160
rect 12238 -14200 12298 -14194
rect -22 -14752 12 -14736
rect 2582 -14244 2616 -14228
rect -7656 -14786 -7596 -14784
rect -6642 -14786 -6582 -14784
rect -2568 -14786 -2508 -14784
rect -1552 -14786 -1492 -14784
rect -8952 -14820 -8936 -14786
rect -8380 -14820 -8364 -14786
rect -7934 -14820 -7918 -14786
rect -7362 -14820 -7346 -14786
rect -6916 -14820 -6900 -14786
rect -6344 -14820 -6328 -14786
rect -5898 -14820 -5882 -14786
rect -5326 -14820 -5310 -14786
rect -4880 -14820 -4864 -14786
rect -4308 -14820 -4292 -14786
rect -3862 -14820 -3846 -14786
rect -3290 -14820 -3274 -14786
rect -2844 -14820 -2828 -14786
rect -2272 -14820 -2256 -14786
rect -1826 -14820 -1810 -14786
rect -1254 -14820 -1238 -14786
rect -808 -14820 -792 -14786
rect -236 -14820 -220 -14786
rect 2582 -14836 2616 -14820
rect 3600 -14244 3634 -14228
rect 3600 -14836 3634 -14820
rect 4618 -14244 4652 -14228
rect 4618 -14836 4652 -14820
rect 5636 -14244 5670 -14228
rect 5636 -14836 5670 -14820
rect 6654 -14244 6688 -14228
rect 6654 -14836 6688 -14820
rect 7672 -14244 7706 -14228
rect 7672 -14836 7706 -14820
rect 8690 -14244 8724 -14228
rect 8690 -14836 8724 -14820
rect 9708 -14244 9742 -14228
rect 9708 -14836 9742 -14820
rect 10726 -14244 10760 -14228
rect 10726 -14836 10760 -14820
rect 11744 -14244 11778 -14228
rect 11744 -14836 11778 -14820
rect 12762 -14244 12796 -14228
rect 12762 -14836 12796 -14820
rect 13780 -14244 13814 -14228
rect 13780 -14836 13814 -14820
rect 14798 -14244 14832 -14228
rect 14798 -14836 14832 -14820
rect 15816 -14244 15850 -14228
rect 15816 -14836 15850 -14820
rect 16834 -14244 16868 -14228
rect 16834 -14836 16868 -14820
rect 17852 -14244 17886 -14228
rect 17852 -14836 17886 -14820
rect 18870 -14244 18904 -14228
rect 18870 -14836 18904 -14820
rect 19888 -14244 19922 -14228
rect 19888 -14836 19922 -14820
rect 20906 -14244 20940 -14228
rect 20906 -14836 20940 -14820
rect 21924 -14244 21958 -14228
rect 21924 -14836 21958 -14820
rect 22942 -14244 22976 -14228
rect 22942 -14836 22976 -14820
rect 8166 -14870 8226 -14864
rect 10202 -14870 10262 -14864
rect 11222 -14870 11282 -14864
rect 16294 -14870 16354 -14864
rect -8952 -14928 -8936 -14894
rect -8380 -14928 -8364 -14894
rect -7934 -14928 -7918 -14894
rect -7362 -14928 -7346 -14894
rect -6916 -14928 -6900 -14894
rect -6344 -14928 -6328 -14894
rect -5898 -14928 -5882 -14894
rect -5326 -14928 -5310 -14894
rect -4880 -14928 -4864 -14894
rect -4308 -14928 -4292 -14894
rect -3862 -14928 -3846 -14894
rect -3290 -14928 -3274 -14894
rect -2844 -14928 -2828 -14894
rect -2272 -14928 -2256 -14894
rect -1826 -14928 -1810 -14894
rect -1254 -14928 -1238 -14894
rect -808 -14928 -792 -14894
rect -236 -14928 -220 -14894
rect 2814 -14904 2830 -14870
rect 3386 -14904 3402 -14870
rect 3832 -14904 3848 -14870
rect 4404 -14904 4420 -14870
rect 4850 -14904 4866 -14870
rect 5422 -14904 5438 -14870
rect 5868 -14904 5884 -14870
rect 6440 -14904 6456 -14870
rect 6886 -14904 6902 -14870
rect 7458 -14904 7474 -14870
rect 7904 -14904 7920 -14870
rect 8476 -14904 8492 -14870
rect 8922 -14904 8938 -14870
rect 9494 -14904 9510 -14870
rect 9940 -14904 9956 -14870
rect 10512 -14904 10528 -14870
rect 10958 -14904 10974 -14870
rect 11530 -14904 11546 -14870
rect 11976 -14904 11992 -14870
rect 12548 -14904 12564 -14870
rect 12994 -14904 13010 -14870
rect 13566 -14904 13582 -14870
rect 14012 -14904 14028 -14870
rect 14584 -14904 14600 -14870
rect 15030 -14904 15046 -14870
rect 15602 -14904 15618 -14870
rect 16048 -14904 16064 -14870
rect 16620 -14904 16636 -14870
rect 17066 -14904 17082 -14870
rect 17638 -14904 17654 -14870
rect 18084 -14904 18100 -14870
rect 18656 -14904 18672 -14870
rect 19102 -14904 19118 -14870
rect 19674 -14904 19690 -14870
rect 20120 -14904 20136 -14870
rect 20692 -14904 20708 -14870
rect 21138 -14904 21154 -14870
rect 21710 -14904 21726 -14870
rect 22156 -14904 22172 -14870
rect 22728 -14904 22744 -14870
rect -9184 -14978 -9150 -14962
rect -9184 -15570 -9150 -15554
rect -8166 -14978 -8132 -14962
rect -8166 -15570 -8132 -15554
rect -7148 -14978 -7114 -14962
rect -7148 -15570 -7114 -15554
rect -6130 -14978 -6096 -14962
rect -6130 -15570 -6096 -15554
rect -5112 -14978 -5078 -14962
rect -5112 -15570 -5078 -15554
rect -4094 -14978 -4060 -14962
rect -4094 -15570 -4060 -15554
rect -3076 -14978 -3042 -14962
rect -3076 -15570 -3042 -15554
rect -2058 -14978 -2024 -14962
rect -2058 -15570 -2024 -15554
rect -1040 -14978 -1006 -14962
rect -1040 -15570 -1006 -15554
rect -22 -14978 12 -14962
rect 2814 -15426 2830 -15392
rect 3386 -15426 3402 -15392
rect 3832 -15426 3848 -15392
rect 4404 -15426 4420 -15392
rect 4850 -15426 4866 -15392
rect 5422 -15426 5438 -15392
rect 5868 -15426 5884 -15392
rect 6440 -15426 6456 -15392
rect 6886 -15426 6902 -15392
rect 7458 -15426 7474 -15392
rect 7904 -15426 7920 -15392
rect 8476 -15426 8492 -15392
rect 8922 -15426 8938 -15392
rect 9494 -15426 9510 -15392
rect 9940 -15426 9956 -15392
rect 10512 -15426 10528 -15392
rect 10958 -15426 10974 -15392
rect 11530 -15426 11546 -15392
rect 11976 -15426 11992 -15392
rect 12548 -15426 12564 -15392
rect 12994 -15426 13010 -15392
rect 13566 -15426 13582 -15392
rect 14012 -15426 14028 -15392
rect 14584 -15426 14600 -15392
rect 15030 -15426 15046 -15392
rect 15602 -15426 15618 -15392
rect 16048 -15426 16064 -15392
rect 16620 -15426 16636 -15392
rect 17066 -15426 17082 -15392
rect 17638 -15426 17654 -15392
rect 18084 -15426 18100 -15392
rect 18656 -15426 18672 -15392
rect 19102 -15426 19118 -15392
rect 19674 -15426 19690 -15392
rect 20120 -15426 20136 -15392
rect 20692 -15426 20708 -15392
rect 21138 -15426 21154 -15392
rect 21710 -15426 21726 -15392
rect 22156 -15426 22172 -15392
rect 22728 -15426 22744 -15392
rect 4100 -15430 4160 -15426
rect 5116 -15430 5176 -15426
rect 9192 -15434 9252 -15426
rect 13258 -15430 13318 -15426
rect 15292 -15430 15352 -15426
rect 21404 -15430 21464 -15426
rect -22 -15570 12 -15554
rect 2582 -15476 2616 -15460
rect -8952 -15638 -8936 -15604
rect -8380 -15638 -8364 -15604
rect -7934 -15638 -7918 -15604
rect -7362 -15638 -7346 -15604
rect -6916 -15638 -6900 -15604
rect -6344 -15638 -6328 -15604
rect -5898 -15638 -5882 -15604
rect -5326 -15638 -5310 -15604
rect -4880 -15638 -4864 -15604
rect -4308 -15638 -4292 -15604
rect -3862 -15638 -3846 -15604
rect -3290 -15638 -3274 -15604
rect -2844 -15638 -2828 -15604
rect -2272 -15638 -2256 -15604
rect -1826 -15638 -1810 -15604
rect -1254 -15638 -1238 -15604
rect -808 -15638 -792 -15604
rect -236 -15638 -220 -15604
rect -8952 -15746 -8936 -15712
rect -8380 -15746 -8364 -15712
rect -7934 -15746 -7918 -15712
rect -7362 -15746 -7346 -15712
rect -6916 -15746 -6900 -15712
rect -6344 -15746 -6328 -15712
rect -5898 -15746 -5882 -15712
rect -5326 -15746 -5310 -15712
rect -4880 -15746 -4864 -15712
rect -4308 -15746 -4292 -15712
rect -3862 -15746 -3846 -15712
rect -3290 -15746 -3274 -15712
rect -2844 -15746 -2828 -15712
rect -2272 -15746 -2256 -15712
rect -1826 -15746 -1810 -15712
rect -1254 -15746 -1238 -15712
rect -808 -15746 -792 -15712
rect -236 -15746 -220 -15712
rect -3596 -15748 -3536 -15746
rect -9184 -15796 -9150 -15780
rect -9184 -16388 -9150 -16372
rect -8166 -15796 -8132 -15780
rect -8166 -16388 -8132 -16372
rect -7148 -15796 -7114 -15780
rect -7148 -16388 -7114 -16372
rect -6130 -15796 -6096 -15780
rect -6130 -16388 -6096 -16372
rect -5112 -15796 -5078 -15780
rect -5112 -16388 -5078 -16372
rect -4094 -15796 -4060 -15780
rect -4094 -16388 -4060 -16372
rect -3076 -15796 -3042 -15780
rect -3076 -16388 -3042 -16372
rect -2058 -15796 -2024 -15780
rect -2058 -16388 -2024 -16372
rect -1040 -15796 -1006 -15780
rect -1040 -16388 -1006 -16372
rect -22 -15796 12 -15780
rect 2582 -16068 2616 -16052
rect 3600 -15476 3634 -15460
rect 3600 -16068 3634 -16052
rect 4618 -15476 4652 -15460
rect 4618 -16068 4652 -16052
rect 5636 -15476 5670 -15460
rect 5636 -16068 5670 -16052
rect 6654 -15476 6688 -15460
rect 6654 -16068 6688 -16052
rect 7672 -15476 7706 -15460
rect 7672 -16068 7706 -16052
rect 8690 -15476 8724 -15460
rect 8690 -16068 8724 -16052
rect 9708 -15476 9742 -15460
rect 9708 -16068 9742 -16052
rect 10726 -15476 10760 -15460
rect 10726 -16068 10760 -16052
rect 11744 -15476 11778 -15460
rect 11744 -16068 11778 -16052
rect 12762 -15476 12796 -15460
rect 12762 -16068 12796 -16052
rect 13780 -15476 13814 -15460
rect 13780 -16068 13814 -16052
rect 14798 -15476 14832 -15460
rect 14798 -16068 14832 -16052
rect 15816 -15476 15850 -15460
rect 15816 -16068 15850 -16052
rect 16834 -15476 16868 -15460
rect 16834 -16068 16868 -16052
rect 17852 -15476 17886 -15460
rect 17852 -16068 17886 -16052
rect 18870 -15476 18904 -15460
rect 18870 -16068 18904 -16052
rect 19888 -15476 19922 -15460
rect 19888 -16068 19922 -16052
rect 20906 -15476 20940 -15460
rect 20906 -16068 20940 -16052
rect 21924 -15476 21958 -15460
rect 21924 -16068 21958 -16052
rect 22942 -15476 22976 -15460
rect 22976 -16052 22982 -16004
rect 22942 -16068 22976 -16052
rect 6126 -16102 6186 -16100
rect 2814 -16136 2830 -16102
rect 3386 -16136 3402 -16102
rect 3832 -16136 3848 -16102
rect 4404 -16136 4420 -16102
rect 4850 -16136 4866 -16102
rect 5422 -16136 5438 -16102
rect 5868 -16136 5884 -16102
rect 6440 -16136 6456 -16102
rect 6886 -16136 6902 -16102
rect 7458 -16136 7474 -16102
rect 7904 -16136 7920 -16102
rect 8476 -16136 8492 -16102
rect 8922 -16136 8938 -16102
rect 9494 -16136 9510 -16102
rect 9940 -16136 9956 -16102
rect 10512 -16136 10528 -16102
rect 10958 -16136 10974 -16102
rect 11530 -16136 11546 -16102
rect 11976 -16136 11992 -16102
rect 12548 -16136 12564 -16102
rect 12994 -16136 13010 -16102
rect 13566 -16136 13582 -16102
rect 14012 -16136 14028 -16102
rect 14584 -16136 14600 -16102
rect 15030 -16136 15046 -16102
rect 15602 -16136 15618 -16102
rect 16048 -16136 16064 -16102
rect 16620 -16136 16636 -16102
rect 17066 -16136 17082 -16102
rect 17638 -16136 17654 -16102
rect 18084 -16136 18100 -16102
rect 18656 -16136 18672 -16102
rect 19102 -16136 19118 -16102
rect 19674 -16136 19690 -16102
rect 20120 -16136 20136 -16102
rect 20692 -16136 20708 -16102
rect 21138 -16136 21154 -16102
rect 21710 -16136 21726 -16102
rect 22156 -16136 22172 -16102
rect 22728 -16136 22744 -16102
rect 8160 -16140 8220 -16136
rect 17318 -16150 17378 -16136
rect 18352 -16150 18412 -16136
rect -22 -16388 12 -16372
rect -7670 -16422 -7610 -16420
rect -6656 -16422 -6596 -16420
rect -2582 -16422 -2522 -16420
rect -1566 -16422 -1506 -16420
rect -8952 -16456 -8936 -16422
rect -8380 -16456 -8364 -16422
rect -7934 -16456 -7918 -16422
rect -7362 -16456 -7346 -16422
rect -6916 -16456 -6900 -16422
rect -6344 -16456 -6328 -16422
rect -5898 -16456 -5882 -16422
rect -5326 -16456 -5310 -16422
rect -4880 -16456 -4864 -16422
rect -4308 -16456 -4292 -16422
rect -3862 -16456 -3846 -16422
rect -3290 -16456 -3274 -16422
rect -2844 -16456 -2828 -16422
rect -2272 -16456 -2256 -16422
rect -1826 -16456 -1810 -16422
rect -1254 -16456 -1238 -16422
rect -808 -16456 -792 -16422
rect -236 -16456 -220 -16422
rect -8952 -16564 -8936 -16530
rect -8380 -16564 -8364 -16530
rect -7934 -16564 -7918 -16530
rect -7362 -16564 -7346 -16530
rect -6916 -16564 -6900 -16530
rect -6344 -16564 -6328 -16530
rect -5898 -16564 -5882 -16530
rect -5326 -16564 -5310 -16530
rect -4880 -16564 -4864 -16530
rect -4308 -16564 -4292 -16530
rect -3862 -16564 -3846 -16530
rect -3290 -16564 -3274 -16530
rect -2844 -16564 -2828 -16530
rect -2272 -16564 -2256 -16530
rect -1826 -16564 -1810 -16530
rect -1254 -16564 -1238 -16530
rect -808 -16564 -792 -16530
rect -236 -16564 -220 -16530
rect -9184 -16614 -9150 -16598
rect -9184 -17206 -9150 -17190
rect -8166 -16614 -8132 -16598
rect -8166 -17206 -8132 -17190
rect -7148 -16614 -7114 -16598
rect -7148 -17206 -7114 -17190
rect -6130 -16614 -6096 -16598
rect -6130 -17206 -6096 -17190
rect -5112 -16614 -5078 -16598
rect -5112 -17206 -5078 -17190
rect -4094 -16614 -4060 -16598
rect -4094 -17206 -4060 -17190
rect -3076 -16614 -3042 -16598
rect -3076 -17206 -3042 -17190
rect -2058 -16614 -2024 -16598
rect -2058 -17206 -2024 -17190
rect -1040 -16614 -1006 -16598
rect -1040 -17206 -1006 -17190
rect -22 -16614 12 -16598
rect 2812 -16660 2828 -16626
rect 3384 -16660 3400 -16626
rect 3830 -16660 3846 -16626
rect 4402 -16660 4418 -16626
rect 4848 -16660 4864 -16626
rect 5420 -16660 5436 -16626
rect 5866 -16660 5882 -16626
rect 6438 -16660 6454 -16626
rect 6884 -16660 6900 -16626
rect 7456 -16660 7472 -16626
rect 7902 -16660 7918 -16626
rect 8474 -16660 8490 -16626
rect 8920 -16660 8936 -16626
rect 9492 -16660 9508 -16626
rect 9938 -16660 9954 -16626
rect 10510 -16660 10526 -16626
rect 10956 -16660 10972 -16626
rect 11528 -16660 11544 -16626
rect 11974 -16660 11990 -16626
rect 12546 -16660 12562 -16626
rect 12992 -16660 13008 -16626
rect 13564 -16660 13580 -16626
rect 14010 -16660 14026 -16626
rect 14582 -16660 14598 -16626
rect 15028 -16660 15044 -16626
rect 15600 -16660 15616 -16626
rect 16046 -16660 16062 -16626
rect 16618 -16660 16634 -16626
rect 17064 -16660 17080 -16626
rect 17636 -16660 17652 -16626
rect 18082 -16660 18098 -16626
rect 18654 -16660 18670 -16626
rect 19100 -16660 19116 -16626
rect 19672 -16660 19688 -16626
rect 20118 -16660 20134 -16626
rect 20690 -16660 20706 -16626
rect 21136 -16660 21152 -16626
rect 21708 -16660 21724 -16626
rect 22154 -16660 22170 -16626
rect 22726 -16660 22742 -16626
rect 5122 -16664 5182 -16660
rect -22 -17206 12 -17190
rect 2580 -16710 2614 -16694
rect -7666 -17240 -7606 -17238
rect -6652 -17240 -6592 -17238
rect -2578 -17240 -2518 -17238
rect -1562 -17240 -1502 -17238
rect -8952 -17274 -8936 -17240
rect -8380 -17274 -8364 -17240
rect -7934 -17274 -7918 -17240
rect -7362 -17274 -7346 -17240
rect -6916 -17274 -6900 -17240
rect -6344 -17274 -6328 -17240
rect -5898 -17274 -5882 -17240
rect -5326 -17274 -5310 -17240
rect -4880 -17274 -4864 -17240
rect -4308 -17274 -4292 -17240
rect -3862 -17274 -3846 -17240
rect -3290 -17274 -3274 -17240
rect -2844 -17274 -2828 -17240
rect -2272 -17274 -2256 -17240
rect -1826 -17274 -1810 -17240
rect -1254 -17274 -1238 -17240
rect -808 -17274 -792 -17240
rect -236 -17274 -220 -17240
rect 2580 -17302 2614 -17286
rect 3598 -16710 3632 -16694
rect 3598 -17302 3632 -17286
rect 4616 -16710 4650 -16694
rect 4616 -17302 4650 -17286
rect 5634 -16710 5668 -16694
rect 5634 -17302 5668 -17286
rect 6652 -16710 6686 -16694
rect 6652 -17302 6686 -17286
rect 7670 -16710 7704 -16694
rect 7670 -17302 7704 -17286
rect 8688 -16710 8722 -16694
rect 8688 -17302 8722 -17286
rect 9706 -16710 9740 -16694
rect 9706 -17302 9740 -17286
rect 10724 -16710 10758 -16694
rect 10724 -17302 10758 -17286
rect 11742 -16710 11776 -16694
rect 11742 -17302 11776 -17286
rect 12760 -16710 12794 -16694
rect 12760 -17302 12794 -17286
rect 13778 -16710 13812 -16694
rect 13778 -17302 13812 -17286
rect 14796 -16710 14830 -16694
rect 14796 -17302 14830 -17286
rect 15814 -16710 15848 -16694
rect 15814 -17302 15848 -17286
rect 16832 -16710 16866 -16694
rect 16832 -17302 16866 -17286
rect 17850 -16710 17884 -16694
rect 17850 -17302 17884 -17286
rect 18868 -16710 18902 -16694
rect 18868 -17302 18902 -17286
rect 19886 -16710 19920 -16694
rect 19886 -17302 19920 -17286
rect 20904 -16710 20938 -16694
rect 20904 -17302 20938 -17286
rect 21922 -16710 21956 -16694
rect 21922 -17302 21956 -17286
rect 22940 -16710 22974 -16694
rect 22940 -17302 22974 -17286
rect 10190 -17336 10250 -17332
rect 11218 -17336 11278 -17334
rect 13262 -17336 13322 -17332
rect -8952 -17382 -8936 -17348
rect -8380 -17382 -8364 -17348
rect -7934 -17382 -7918 -17348
rect -7362 -17382 -7346 -17348
rect -6916 -17382 -6900 -17348
rect -6344 -17382 -6328 -17348
rect -5898 -17382 -5882 -17348
rect -5326 -17382 -5310 -17348
rect -4880 -17382 -4864 -17348
rect -4308 -17382 -4292 -17348
rect -3862 -17382 -3846 -17348
rect -3290 -17382 -3274 -17348
rect -2844 -17382 -2828 -17348
rect -2272 -17382 -2256 -17348
rect -1826 -17382 -1810 -17348
rect -1254 -17382 -1238 -17348
rect -808 -17382 -792 -17348
rect -236 -17382 -220 -17348
rect 2812 -17370 2828 -17336
rect 3384 -17370 3400 -17336
rect 3830 -17370 3846 -17336
rect 4402 -17370 4418 -17336
rect 4848 -17370 4864 -17336
rect 5420 -17370 5436 -17336
rect 5866 -17370 5882 -17336
rect 6438 -17370 6454 -17336
rect 6884 -17370 6900 -17336
rect 7456 -17370 7472 -17336
rect 7902 -17370 7918 -17336
rect 8474 -17370 8490 -17336
rect 8920 -17370 8936 -17336
rect 9492 -17370 9508 -17336
rect 9938 -17370 9954 -17336
rect 10510 -17370 10526 -17336
rect 10956 -17370 10972 -17336
rect 11528 -17370 11544 -17336
rect 11974 -17370 11990 -17336
rect 12546 -17370 12562 -17336
rect 12992 -17370 13008 -17336
rect 13564 -17370 13580 -17336
rect 14010 -17370 14026 -17336
rect 14582 -17370 14598 -17336
rect 15028 -17370 15044 -17336
rect 15600 -17370 15616 -17336
rect 16046 -17370 16062 -17336
rect 16618 -17370 16634 -17336
rect 17064 -17370 17080 -17336
rect 17636 -17370 17652 -17336
rect 18082 -17370 18098 -17336
rect 18654 -17370 18670 -17336
rect 19100 -17370 19116 -17336
rect 19672 -17370 19688 -17336
rect 20118 -17370 20134 -17336
rect 20690 -17370 20706 -17336
rect 21136 -17370 21152 -17336
rect 21708 -17370 21724 -17336
rect 22154 -17370 22170 -17336
rect 22726 -17370 22742 -17336
rect -9184 -17432 -9150 -17416
rect -9184 -18024 -9150 -18008
rect -8166 -17432 -8132 -17416
rect -8166 -18024 -8132 -18008
rect -7148 -17432 -7114 -17416
rect -7148 -18024 -7114 -18008
rect -6130 -17432 -6096 -17416
rect -6130 -18024 -6096 -18008
rect -5112 -17432 -5078 -17416
rect -5112 -18024 -5078 -18008
rect -4094 -17432 -4060 -17416
rect -4094 -18024 -4060 -18008
rect -3076 -17432 -3042 -17416
rect -3076 -18024 -3042 -18008
rect -2058 -17432 -2024 -17416
rect -2058 -18024 -2024 -18008
rect -1040 -17432 -1006 -17416
rect -1040 -18024 -1006 -18008
rect -22 -17432 12 -17416
rect 2812 -17894 2828 -17860
rect 3384 -17894 3400 -17860
rect 3830 -17894 3846 -17860
rect 4402 -17894 4418 -17860
rect 4848 -17894 4864 -17860
rect 5420 -17894 5436 -17860
rect 5866 -17894 5882 -17860
rect 6438 -17894 6454 -17860
rect 6884 -17894 6900 -17860
rect 7456 -17894 7472 -17860
rect 7902 -17894 7918 -17860
rect 8474 -17894 8490 -17860
rect 8920 -17894 8936 -17860
rect 9492 -17894 9508 -17860
rect 9938 -17894 9954 -17860
rect 10510 -17894 10526 -17860
rect 10956 -17894 10972 -17860
rect 11528 -17894 11544 -17860
rect 11974 -17894 11990 -17860
rect 12546 -17894 12562 -17860
rect 12992 -17894 13008 -17860
rect 13564 -17894 13580 -17860
rect 14010 -17894 14026 -17860
rect 14582 -17894 14598 -17860
rect 15028 -17894 15044 -17860
rect 15600 -17894 15616 -17860
rect 16046 -17894 16062 -17860
rect 16618 -17894 16634 -17860
rect 17064 -17894 17080 -17860
rect 17636 -17894 17652 -17860
rect 18082 -17894 18098 -17860
rect 18654 -17894 18670 -17860
rect 19100 -17894 19116 -17860
rect 19672 -17894 19688 -17860
rect 20118 -17894 20134 -17860
rect 20690 -17894 20706 -17860
rect 21136 -17894 21152 -17860
rect 21708 -17894 21724 -17860
rect 22154 -17894 22170 -17860
rect 22726 -17894 22742 -17860
rect -22 -18024 12 -18008
rect 2580 -17944 2614 -17928
rect -8692 -18058 -8632 -18056
rect -7666 -18058 -7606 -18054
rect -6652 -18058 -6592 -18054
rect -5632 -18058 -5572 -18056
rect -4610 -18058 -4550 -18056
rect -2578 -18058 -2518 -18054
rect -1562 -18058 -1502 -18054
rect -542 -18058 -482 -18056
rect -8952 -18092 -8936 -18058
rect -8380 -18092 -8364 -18058
rect -7934 -18092 -7918 -18058
rect -7362 -18092 -7346 -18058
rect -6916 -18092 -6900 -18058
rect -6344 -18092 -6328 -18058
rect -5898 -18092 -5882 -18058
rect -5326 -18092 -5310 -18058
rect -4880 -18092 -4864 -18058
rect -4308 -18092 -4292 -18058
rect -3862 -18092 -3846 -18058
rect -3290 -18092 -3274 -18058
rect -2844 -18092 -2828 -18058
rect -2272 -18092 -2256 -18058
rect -1826 -18092 -1810 -18058
rect -1254 -18092 -1238 -18058
rect -808 -18092 -792 -18058
rect -236 -18092 -220 -18058
rect -8952 -18200 -8936 -18166
rect -8380 -18200 -8364 -18166
rect -7934 -18200 -7918 -18166
rect -7362 -18200 -7346 -18166
rect -6916 -18200 -6900 -18166
rect -6344 -18200 -6328 -18166
rect -5898 -18200 -5882 -18166
rect -5326 -18200 -5310 -18166
rect -4880 -18200 -4864 -18166
rect -4308 -18200 -4292 -18166
rect -3862 -18200 -3846 -18166
rect -3290 -18200 -3274 -18166
rect -2844 -18200 -2828 -18166
rect -2272 -18200 -2256 -18166
rect -1826 -18200 -1810 -18166
rect -1254 -18200 -1238 -18166
rect -808 -18200 -792 -18166
rect -236 -18200 -220 -18166
rect -9184 -18250 -9150 -18234
rect -9184 -18842 -9150 -18826
rect -8166 -18250 -8132 -18234
rect -8166 -18842 -8132 -18826
rect -7148 -18250 -7114 -18234
rect -7148 -18842 -7114 -18826
rect -6130 -18250 -6096 -18234
rect -6130 -18842 -6096 -18826
rect -5112 -18250 -5078 -18234
rect -5112 -18842 -5078 -18826
rect -4094 -18250 -4060 -18234
rect -4094 -18842 -4060 -18826
rect -3076 -18250 -3042 -18234
rect -3076 -18842 -3042 -18826
rect -2058 -18250 -2024 -18234
rect -2058 -18842 -2024 -18826
rect -1040 -18250 -1006 -18234
rect -1040 -18842 -1006 -18826
rect -22 -18250 12 -18234
rect 2580 -18536 2614 -18520
rect 3598 -17944 3632 -17928
rect 3598 -18536 3632 -18520
rect 4616 -17944 4650 -17928
rect 4616 -18536 4650 -18520
rect 5634 -17944 5668 -17928
rect 5634 -18536 5668 -18520
rect 6652 -17944 6686 -17928
rect 6652 -18536 6686 -18520
rect 7670 -17944 7704 -17928
rect 7670 -18536 7704 -18520
rect 8688 -17944 8722 -17928
rect 8688 -18536 8722 -18520
rect 9706 -17944 9740 -17928
rect 9706 -18536 9740 -18520
rect 10724 -17944 10758 -17928
rect 10724 -18536 10758 -18520
rect 11742 -17944 11776 -17928
rect 11742 -18536 11776 -18520
rect 12760 -17944 12794 -17928
rect 12760 -18536 12794 -18520
rect 13778 -17944 13812 -17928
rect 13778 -18536 13812 -18520
rect 14796 -17944 14830 -17928
rect 14796 -18536 14830 -18520
rect 15814 -17944 15848 -17928
rect 15814 -18536 15848 -18520
rect 16832 -17944 16866 -17928
rect 16832 -18536 16866 -18520
rect 17850 -17944 17884 -17928
rect 17850 -18536 17884 -18520
rect 18868 -17944 18902 -17928
rect 18868 -18536 18902 -18520
rect 19886 -17944 19920 -17928
rect 19886 -18536 19920 -18520
rect 20904 -17944 20938 -17928
rect 20904 -18536 20938 -18520
rect 21922 -17944 21956 -17928
rect 21922 -18536 21956 -18520
rect 22940 -17944 22974 -17928
rect 22940 -18536 22974 -18520
rect 2812 -18604 2828 -18570
rect 3384 -18604 3400 -18570
rect 3830 -18604 3846 -18570
rect 4402 -18604 4418 -18570
rect 4848 -18604 4864 -18570
rect 5420 -18604 5436 -18570
rect 5866 -18604 5882 -18570
rect 6438 -18604 6454 -18570
rect 6884 -18604 6900 -18570
rect 7456 -18604 7472 -18570
rect 7902 -18604 7918 -18570
rect 8474 -18604 8490 -18570
rect 8920 -18604 8936 -18570
rect 9492 -18604 9508 -18570
rect 9938 -18604 9954 -18570
rect 10510 -18604 10526 -18570
rect 10956 -18604 10972 -18570
rect 11528 -18604 11544 -18570
rect 11974 -18604 11990 -18570
rect 12546 -18604 12562 -18570
rect 12992 -18604 13008 -18570
rect 13564 -18604 13580 -18570
rect 14010 -18604 14026 -18570
rect 14582 -18604 14598 -18570
rect 15028 -18604 15044 -18570
rect 15600 -18604 15616 -18570
rect 16046 -18604 16062 -18570
rect 16618 -18604 16634 -18570
rect 17064 -18604 17080 -18570
rect 17636 -18604 17652 -18570
rect 18082 -18604 18098 -18570
rect 18654 -18604 18670 -18570
rect 19100 -18604 19116 -18570
rect 19672 -18604 19688 -18570
rect 20118 -18604 20134 -18570
rect 20690 -18604 20706 -18570
rect 21136 -18604 21152 -18570
rect 21708 -18604 21724 -18570
rect 22154 -18604 22170 -18570
rect 22726 -18604 22742 -18570
rect -22 -18842 12 -18826
rect -8952 -18910 -8936 -18876
rect -8380 -18910 -8364 -18876
rect -7934 -18910 -7918 -18876
rect -7362 -18910 -7346 -18876
rect -6916 -18910 -6900 -18876
rect -6344 -18910 -6328 -18876
rect -5898 -18910 -5882 -18876
rect -5326 -18910 -5310 -18876
rect -4880 -18910 -4864 -18876
rect -4308 -18910 -4292 -18876
rect -3862 -18910 -3846 -18876
rect -3290 -18910 -3274 -18876
rect -2844 -18910 -2828 -18876
rect -2272 -18910 -2256 -18876
rect -1826 -18910 -1810 -18876
rect -1254 -18910 -1238 -18876
rect -808 -18910 -792 -18876
rect -236 -18910 -220 -18876
rect 2812 -19126 2828 -19092
rect 3384 -19126 3400 -19092
rect 3830 -19126 3846 -19092
rect 4402 -19126 4418 -19092
rect 4848 -19126 4864 -19092
rect 5420 -19126 5436 -19092
rect 5866 -19126 5882 -19092
rect 6438 -19126 6454 -19092
rect 6884 -19126 6900 -19092
rect 7456 -19126 7472 -19092
rect 7902 -19126 7918 -19092
rect 8474 -19126 8490 -19092
rect 8920 -19126 8936 -19092
rect 9492 -19126 9508 -19092
rect 9938 -19126 9954 -19092
rect 10510 -19126 10526 -19092
rect 10956 -19126 10972 -19092
rect 11528 -19126 11544 -19092
rect 11974 -19126 11990 -19092
rect 12546 -19126 12562 -19092
rect 12992 -19126 13008 -19092
rect 13564 -19126 13580 -19092
rect 14010 -19126 14026 -19092
rect 14582 -19126 14598 -19092
rect 15028 -19126 15044 -19092
rect 15600 -19126 15616 -19092
rect 16046 -19126 16062 -19092
rect 16618 -19126 16634 -19092
rect 17064 -19126 17080 -19092
rect 17636 -19126 17652 -19092
rect 18082 -19126 18098 -19092
rect 18654 -19126 18670 -19092
rect 19100 -19126 19116 -19092
rect 19672 -19126 19688 -19092
rect 20118 -19126 20134 -19092
rect 20690 -19126 20706 -19092
rect 21136 -19126 21152 -19092
rect 21708 -19126 21724 -19092
rect 22154 -19126 22170 -19092
rect 22726 -19126 22742 -19092
rect 2580 -19176 2614 -19160
rect 2580 -19768 2614 -19752
rect 3598 -19176 3632 -19160
rect 3598 -19768 3632 -19752
rect 4616 -19176 4650 -19160
rect 4616 -19768 4650 -19752
rect 5634 -19176 5668 -19160
rect 5634 -19768 5668 -19752
rect 6652 -19176 6686 -19160
rect 6652 -19768 6686 -19752
rect 7670 -19176 7704 -19160
rect 7670 -19768 7704 -19752
rect 8688 -19176 8722 -19160
rect 8688 -19768 8722 -19752
rect 9706 -19176 9740 -19160
rect 9706 -19768 9740 -19752
rect 10724 -19176 10758 -19160
rect 10724 -19768 10758 -19752
rect 11742 -19176 11776 -19160
rect 11742 -19768 11776 -19752
rect 12760 -19176 12794 -19160
rect 12760 -19768 12794 -19752
rect 13778 -19176 13812 -19160
rect 13778 -19768 13812 -19752
rect 14796 -19176 14830 -19160
rect 14796 -19768 14830 -19752
rect 15814 -19176 15848 -19160
rect 15814 -19768 15848 -19752
rect 16832 -19176 16866 -19160
rect 16832 -19768 16866 -19752
rect 17850 -19176 17884 -19160
rect 17850 -19768 17884 -19752
rect 18868 -19176 18902 -19160
rect 18868 -19768 18902 -19752
rect 19886 -19176 19920 -19160
rect 19886 -19768 19920 -19752
rect 20904 -19176 20938 -19160
rect 20904 -19768 20938 -19752
rect 21922 -19176 21956 -19160
rect 21922 -19768 21956 -19752
rect 22940 -19176 22974 -19160
rect 22940 -19768 22974 -19752
rect 11230 -19802 11290 -19800
rect 13274 -19802 13334 -19798
rect 21408 -19802 21468 -19800
rect 2812 -19836 2828 -19802
rect 3384 -19836 3400 -19802
rect 3830 -19836 3846 -19802
rect 4402 -19836 4418 -19802
rect 4848 -19836 4864 -19802
rect 5420 -19836 5436 -19802
rect 5866 -19836 5882 -19802
rect 6438 -19836 6454 -19802
rect 6884 -19836 6900 -19802
rect 7456 -19836 7472 -19802
rect 7902 -19836 7918 -19802
rect 8474 -19836 8490 -19802
rect 8920 -19836 8936 -19802
rect 9492 -19836 9508 -19802
rect 9938 -19836 9954 -19802
rect 10510 -19836 10526 -19802
rect 10956 -19836 10972 -19802
rect 11528 -19836 11544 -19802
rect 11974 -19836 11990 -19802
rect 12546 -19836 12562 -19802
rect 12992 -19836 13008 -19802
rect 13564 -19836 13580 -19802
rect 14010 -19836 14026 -19802
rect 14582 -19836 14598 -19802
rect 15028 -19836 15044 -19802
rect 15600 -19836 15616 -19802
rect 16046 -19836 16062 -19802
rect 16618 -19836 16634 -19802
rect 17064 -19836 17080 -19802
rect 17636 -19836 17652 -19802
rect 18082 -19836 18098 -19802
rect 18654 -19836 18670 -19802
rect 19100 -19836 19116 -19802
rect 19672 -19836 19688 -19802
rect 20118 -19836 20134 -19802
rect 20690 -19836 20706 -19802
rect 21136 -19836 21152 -19802
rect 21708 -19836 21724 -19802
rect 22154 -19836 22170 -19802
rect 22726 -19836 22742 -19802
rect 2812 -20360 2828 -20326
rect 3384 -20360 3400 -20326
rect 3830 -20360 3846 -20326
rect 4402 -20360 4418 -20326
rect 4848 -20360 4864 -20326
rect 5420 -20360 5436 -20326
rect 5866 -20360 5882 -20326
rect 6438 -20360 6454 -20326
rect 6884 -20360 6900 -20326
rect 7456 -20360 7472 -20326
rect 7902 -20360 7918 -20326
rect 8474 -20360 8490 -20326
rect 8920 -20360 8936 -20326
rect 9492 -20360 9508 -20326
rect 9938 -20360 9954 -20326
rect 10510 -20360 10526 -20326
rect 10956 -20360 10972 -20326
rect 11528 -20360 11544 -20326
rect 11974 -20360 11990 -20326
rect 12546 -20360 12562 -20326
rect 12992 -20360 13008 -20326
rect 13564 -20360 13580 -20326
rect 14010 -20360 14026 -20326
rect 14582 -20360 14598 -20326
rect 15028 -20360 15044 -20326
rect 15600 -20360 15616 -20326
rect 16046 -20360 16062 -20326
rect 16618 -20360 16634 -20326
rect 17064 -20360 17080 -20326
rect 17636 -20360 17652 -20326
rect 18082 -20360 18098 -20326
rect 18654 -20360 18670 -20326
rect 19100 -20360 19116 -20326
rect 19672 -20360 19688 -20326
rect 20118 -20360 20134 -20326
rect 20690 -20360 20706 -20326
rect 21136 -20360 21152 -20326
rect 21708 -20360 21724 -20326
rect 22154 -20360 22170 -20326
rect 22726 -20360 22742 -20326
rect 2580 -20410 2614 -20394
rect 2580 -21002 2614 -20986
rect 3598 -20410 3632 -20394
rect 3598 -21002 3632 -20986
rect 4616 -20410 4650 -20394
rect 4616 -21002 4650 -20986
rect 5634 -20410 5668 -20394
rect 5634 -21002 5668 -20986
rect 6652 -20410 6686 -20394
rect 6652 -21002 6686 -20986
rect 7670 -20410 7704 -20394
rect 7670 -21002 7704 -20986
rect 8688 -20410 8722 -20394
rect 8688 -21002 8722 -20986
rect 9706 -20410 9740 -20394
rect 9706 -21002 9740 -20986
rect 10724 -20410 10758 -20394
rect 10724 -21002 10758 -20986
rect 11742 -20410 11776 -20394
rect 11742 -21002 11776 -20986
rect 12760 -20410 12794 -20394
rect 12760 -21002 12794 -20986
rect 13778 -20410 13812 -20394
rect 13778 -21002 13812 -20986
rect 14796 -20410 14830 -20394
rect 14796 -21002 14830 -20986
rect 15814 -20410 15848 -20394
rect 15814 -21002 15848 -20986
rect 16832 -20410 16866 -20394
rect 16832 -21002 16866 -20986
rect 17850 -20410 17884 -20394
rect 17850 -21002 17884 -20986
rect 18868 -20410 18902 -20394
rect 18868 -21002 18902 -20986
rect 19886 -20410 19920 -20394
rect 19886 -21002 19920 -20986
rect 20904 -20410 20938 -20394
rect 20904 -21002 20938 -20986
rect 21922 -20410 21956 -20394
rect 21922 -21002 21956 -20986
rect 22940 -20410 22974 -20394
rect 22940 -21002 22974 -20986
rect 5106 -21036 5166 -21032
rect 2812 -21070 2828 -21036
rect 3384 -21070 3400 -21036
rect 3830 -21070 3846 -21036
rect 4402 -21070 4418 -21036
rect 4848 -21070 4864 -21036
rect 5420 -21070 5436 -21036
rect 5866 -21070 5882 -21036
rect 6438 -21070 6454 -21036
rect 6884 -21070 6900 -21036
rect 7456 -21070 7472 -21036
rect 7902 -21070 7918 -21036
rect 8474 -21070 8490 -21036
rect 8920 -21070 8936 -21036
rect 9492 -21070 9508 -21036
rect 9938 -21070 9954 -21036
rect 10510 -21070 10526 -21036
rect 10956 -21070 10972 -21036
rect 11528 -21070 11544 -21036
rect 11974 -21070 11990 -21036
rect 12546 -21070 12562 -21036
rect 12992 -21070 13008 -21036
rect 13564 -21070 13580 -21036
rect 14010 -21070 14026 -21036
rect 14582 -21070 14598 -21036
rect 15028 -21070 15044 -21036
rect 15600 -21070 15616 -21036
rect 16046 -21070 16062 -21036
rect 16618 -21070 16634 -21036
rect 17064 -21070 17080 -21036
rect 17636 -21070 17652 -21036
rect 18082 -21070 18098 -21036
rect 18654 -21070 18670 -21036
rect 19100 -21070 19116 -21036
rect 19672 -21070 19688 -21036
rect 20118 -21070 20134 -21036
rect 20690 -21070 20706 -21036
rect 21136 -21070 21152 -21036
rect 21708 -21070 21724 -21036
rect 22154 -21070 22170 -21036
rect 22726 -21070 22742 -21036
rect 2812 -21594 2828 -21560
rect 3384 -21594 3400 -21560
rect 3830 -21594 3846 -21560
rect 4402 -21594 4418 -21560
rect 4848 -21594 4864 -21560
rect 5420 -21594 5436 -21560
rect 5866 -21594 5882 -21560
rect 6438 -21594 6454 -21560
rect 6884 -21594 6900 -21560
rect 7456 -21594 7472 -21560
rect 7902 -21594 7918 -21560
rect 8474 -21594 8490 -21560
rect 8920 -21594 8936 -21560
rect 9492 -21594 9508 -21560
rect 9938 -21594 9954 -21560
rect 10510 -21594 10526 -21560
rect 10956 -21594 10972 -21560
rect 11528 -21594 11544 -21560
rect 11974 -21594 11990 -21560
rect 12546 -21594 12562 -21560
rect 12992 -21594 13008 -21560
rect 13564 -21594 13580 -21560
rect 14010 -21594 14026 -21560
rect 14582 -21594 14598 -21560
rect 15028 -21594 15044 -21560
rect 15600 -21594 15616 -21560
rect 16046 -21594 16062 -21560
rect 16618 -21594 16634 -21560
rect 17064 -21594 17080 -21560
rect 17636 -21594 17652 -21560
rect 18082 -21594 18098 -21560
rect 18654 -21594 18670 -21560
rect 19100 -21594 19116 -21560
rect 19672 -21594 19688 -21560
rect 20118 -21594 20134 -21560
rect 20690 -21594 20706 -21560
rect 21136 -21594 21152 -21560
rect 21708 -21594 21724 -21560
rect 22154 -21594 22170 -21560
rect 22726 -21594 22742 -21560
rect 2580 -21644 2614 -21628
rect 2580 -22236 2614 -22220
rect 3598 -21644 3632 -21628
rect 3598 -22236 3632 -22220
rect 4616 -21644 4650 -21628
rect 4616 -22236 4650 -22220
rect 5634 -21644 5668 -21628
rect 5634 -22236 5668 -22220
rect 6652 -21644 6686 -21628
rect 6652 -22236 6686 -22220
rect 7670 -21644 7704 -21628
rect 7670 -22236 7704 -22220
rect 8688 -21644 8722 -21628
rect 8688 -22236 8722 -22220
rect 9706 -21644 9740 -21628
rect 9706 -22236 9740 -22220
rect 10724 -21644 10758 -21628
rect 10724 -22236 10758 -22220
rect 11742 -21644 11776 -21628
rect 11742 -22236 11776 -22220
rect 12760 -21644 12794 -21628
rect 12760 -22236 12794 -22220
rect 13778 -21644 13812 -21628
rect 13778 -22236 13812 -22220
rect 14796 -21644 14830 -21628
rect 14796 -22236 14830 -22220
rect 15814 -21644 15848 -21628
rect 15814 -22236 15848 -22220
rect 16832 -21644 16866 -21628
rect 16832 -22236 16866 -22220
rect 17850 -21644 17884 -21628
rect 17850 -22236 17884 -22220
rect 18868 -21644 18902 -21628
rect 18868 -22236 18902 -22220
rect 19886 -21644 19920 -21628
rect 19886 -22236 19920 -22220
rect 20904 -21644 20938 -21628
rect 20904 -22236 20938 -22220
rect 21922 -21644 21956 -21628
rect 21922 -22236 21956 -22220
rect 22940 -21644 22974 -21628
rect 22940 -22236 22974 -22220
rect 11230 -22270 11290 -22268
rect 13274 -22270 13334 -22266
rect 16312 -22270 16372 -22266
rect 2812 -22304 2828 -22270
rect 3384 -22304 3400 -22270
rect 3830 -22304 3846 -22270
rect 4402 -22304 4418 -22270
rect 4848 -22304 4864 -22270
rect 5420 -22304 5436 -22270
rect 5866 -22304 5882 -22270
rect 6438 -22304 6454 -22270
rect 6884 -22304 6900 -22270
rect 7456 -22304 7472 -22270
rect 7902 -22304 7918 -22270
rect 8474 -22304 8490 -22270
rect 8920 -22304 8936 -22270
rect 9492 -22304 9508 -22270
rect 9938 -22304 9954 -22270
rect 10510 -22304 10526 -22270
rect 10956 -22304 10972 -22270
rect 11528 -22304 11544 -22270
rect 11974 -22304 11990 -22270
rect 12546 -22304 12562 -22270
rect 12992 -22304 13008 -22270
rect 13564 -22304 13580 -22270
rect 14010 -22304 14026 -22270
rect 14582 -22304 14598 -22270
rect 15028 -22304 15044 -22270
rect 15600 -22304 15616 -22270
rect 16046 -22304 16062 -22270
rect 16618 -22304 16634 -22270
rect 17064 -22304 17080 -22270
rect 17636 -22304 17652 -22270
rect 18082 -22304 18098 -22270
rect 18654 -22304 18670 -22270
rect 19100 -22304 19116 -22270
rect 19672 -22304 19688 -22270
rect 20118 -22304 20134 -22270
rect 20690 -22304 20706 -22270
rect 21136 -22304 21152 -22270
rect 21708 -22304 21724 -22270
rect 22154 -22304 22170 -22270
rect 22726 -22304 22742 -22270
rect 2812 -22826 2828 -22792
rect 3384 -22826 3400 -22792
rect 3830 -22826 3846 -22792
rect 4402 -22826 4418 -22792
rect 4848 -22826 4864 -22792
rect 5420 -22826 5436 -22792
rect 5866 -22826 5882 -22792
rect 6438 -22826 6454 -22792
rect 6884 -22826 6900 -22792
rect 7456 -22826 7472 -22792
rect 7902 -22826 7918 -22792
rect 8474 -22826 8490 -22792
rect 8920 -22826 8936 -22792
rect 9492 -22826 9508 -22792
rect 9938 -22826 9954 -22792
rect 10510 -22826 10526 -22792
rect 10956 -22826 10972 -22792
rect 11528 -22826 11544 -22792
rect 11974 -22826 11990 -22792
rect 12546 -22826 12562 -22792
rect 12992 -22826 13008 -22792
rect 13564 -22826 13580 -22792
rect 14010 -22826 14026 -22792
rect 14582 -22826 14598 -22792
rect 15028 -22826 15044 -22792
rect 15600 -22826 15616 -22792
rect 16046 -22826 16062 -22792
rect 16618 -22826 16634 -22792
rect 17064 -22826 17080 -22792
rect 17636 -22826 17652 -22792
rect 18082 -22826 18098 -22792
rect 18654 -22826 18670 -22792
rect 19100 -22826 19116 -22792
rect 19672 -22826 19688 -22792
rect 20118 -22826 20134 -22792
rect 20690 -22826 20706 -22792
rect 21136 -22826 21152 -22792
rect 21708 -22826 21724 -22792
rect 22154 -22826 22170 -22792
rect 22726 -22826 22742 -22792
rect 6134 -22828 6194 -22826
rect 2580 -22876 2614 -22860
rect 2580 -23468 2614 -23452
rect 3598 -22876 3632 -22860
rect 3598 -23468 3632 -23452
rect 4616 -22876 4650 -22860
rect 4616 -23468 4650 -23452
rect 5634 -22876 5668 -22860
rect 5634 -23468 5668 -23452
rect 6652 -22876 6686 -22860
rect 6652 -23468 6686 -23452
rect 7670 -22876 7704 -22860
rect 7670 -23468 7704 -23452
rect 8688 -22876 8722 -22860
rect 8688 -23468 8722 -23452
rect 9706 -22876 9740 -22860
rect 9706 -23468 9740 -23452
rect 10724 -22876 10758 -22860
rect 10724 -23468 10758 -23452
rect 11742 -22876 11776 -22860
rect 11742 -23468 11776 -23452
rect 12760 -22876 12794 -22860
rect 12760 -23468 12794 -23452
rect 13778 -22876 13812 -22860
rect 13778 -23468 13812 -23452
rect 14796 -22876 14830 -22860
rect 14796 -23468 14830 -23452
rect 15814 -22876 15848 -22860
rect 15814 -23468 15848 -23452
rect 16832 -22876 16866 -22860
rect 16832 -23468 16866 -23452
rect 17850 -22876 17884 -22860
rect 17850 -23468 17884 -23452
rect 18868 -22876 18902 -22860
rect 18868 -23468 18902 -23452
rect 19886 -22876 19920 -22860
rect 19886 -23468 19920 -23452
rect 20904 -22876 20938 -22860
rect 21922 -22876 21956 -22860
rect 22940 -22876 22974 -22860
rect 20904 -23468 20938 -23452
rect 22940 -23468 22974 -23452
rect 10206 -23502 10266 -23492
rect 2812 -23536 2828 -23502
rect 3384 -23536 3400 -23502
rect 3830 -23536 3846 -23502
rect 4402 -23536 4418 -23502
rect 4848 -23536 4864 -23502
rect 5420 -23536 5436 -23502
rect 5866 -23536 5882 -23502
rect 6438 -23536 6454 -23502
rect 6884 -23536 6900 -23502
rect 7456 -23536 7472 -23502
rect 7902 -23536 7918 -23502
rect 8474 -23536 8490 -23502
rect 8920 -23536 8936 -23502
rect 9492 -23536 9508 -23502
rect 9938 -23536 9954 -23502
rect 10510 -23536 10526 -23502
rect 10956 -23536 10972 -23502
rect 11528 -23536 11544 -23502
rect 11974 -23536 11990 -23502
rect 12546 -23536 12562 -23502
rect 12992 -23536 13008 -23502
rect 13564 -23536 13580 -23502
rect 14010 -23536 14026 -23502
rect 14582 -23536 14598 -23502
rect 15028 -23536 15044 -23502
rect 15600 -23536 15616 -23502
rect 16046 -23536 16062 -23502
rect 16618 -23536 16634 -23502
rect 17064 -23536 17080 -23502
rect 17636 -23536 17652 -23502
rect 18082 -23536 18098 -23502
rect 18654 -23536 18670 -23502
rect 19100 -23536 19116 -23502
rect 19672 -23536 19688 -23502
rect 20118 -23536 20134 -23502
rect 20690 -23536 20706 -23502
rect 21136 -23536 21152 -23502
rect 21708 -23536 21724 -23502
rect 22154 -23536 22170 -23502
rect 22726 -23536 22742 -23502
rect 2812 -24060 2828 -24026
rect 3384 -24060 3400 -24026
rect 3830 -24060 3846 -24026
rect 4402 -24060 4418 -24026
rect 4848 -24060 4864 -24026
rect 5420 -24060 5436 -24026
rect 5866 -24060 5882 -24026
rect 6438 -24060 6454 -24026
rect 6884 -24060 6900 -24026
rect 7456 -24060 7472 -24026
rect 7902 -24060 7918 -24026
rect 8474 -24060 8490 -24026
rect 8920 -24060 8936 -24026
rect 9492 -24060 9508 -24026
rect 9938 -24060 9954 -24026
rect 10510 -24060 10526 -24026
rect 10956 -24060 10972 -24026
rect 11528 -24060 11544 -24026
rect 11974 -24060 11990 -24026
rect 12546 -24060 12562 -24026
rect 12992 -24060 13008 -24026
rect 13564 -24060 13580 -24026
rect 14010 -24060 14026 -24026
rect 14582 -24060 14598 -24026
rect 15028 -24060 15044 -24026
rect 15600 -24060 15616 -24026
rect 16046 -24060 16062 -24026
rect 16618 -24060 16634 -24026
rect 17064 -24060 17080 -24026
rect 17636 -24060 17652 -24026
rect 18082 -24060 18098 -24026
rect 18654 -24060 18670 -24026
rect 19100 -24060 19116 -24026
rect 19672 -24060 19688 -24026
rect 20118 -24060 20134 -24026
rect 20690 -24060 20706 -24026
rect 21136 -24060 21152 -24026
rect 21708 -24060 21724 -24026
rect 22154 -24060 22170 -24026
rect 22726 -24060 22742 -24026
rect 6120 -24062 6180 -24060
rect 2580 -24110 2614 -24094
rect 2580 -24702 2614 -24686
rect 3598 -24110 3632 -24094
rect 3598 -24702 3632 -24686
rect 4616 -24110 4650 -24094
rect 4616 -24702 4650 -24686
rect 5634 -24110 5668 -24094
rect 5634 -24702 5668 -24686
rect 6652 -24110 6686 -24094
rect 6652 -24702 6686 -24686
rect 7670 -24110 7704 -24094
rect 7670 -24702 7704 -24686
rect 8688 -24110 8722 -24094
rect 8688 -24702 8722 -24686
rect 9706 -24110 9740 -24094
rect 9706 -24702 9740 -24686
rect 10724 -24110 10758 -24094
rect 10724 -24702 10758 -24686
rect 11742 -24110 11776 -24094
rect 11742 -24702 11776 -24686
rect 12760 -24110 12794 -24094
rect 12760 -24702 12794 -24686
rect 13778 -24110 13812 -24094
rect 13778 -24702 13812 -24686
rect 14796 -24110 14830 -24094
rect 14796 -24702 14830 -24686
rect 15814 -24110 15848 -24094
rect 15814 -24702 15848 -24686
rect 16832 -24110 16866 -24094
rect 16832 -24702 16866 -24686
rect 17850 -24110 17884 -24094
rect 17850 -24702 17884 -24686
rect 18868 -24110 18902 -24094
rect 18868 -24702 18902 -24686
rect 19886 -24110 19920 -24094
rect 19886 -24702 19920 -24686
rect 20904 -24110 20938 -24094
rect 20904 -24702 20938 -24686
rect 21922 -24110 21956 -24094
rect 21922 -24702 21956 -24686
rect 22940 -24110 22974 -24094
rect 22940 -24702 22974 -24686
rect 4088 -24736 4148 -24734
rect 10200 -24736 10260 -24734
rect 12234 -24736 12294 -24734
rect 16300 -24736 16360 -24730
rect 20376 -24736 20436 -24734
rect 21392 -24736 21452 -24734
rect 2812 -24770 2828 -24736
rect 3384 -24770 3400 -24736
rect 3830 -24770 3846 -24736
rect 4402 -24770 4418 -24736
rect 4848 -24770 4864 -24736
rect 5420 -24770 5436 -24736
rect 5866 -24770 5882 -24736
rect 6438 -24770 6454 -24736
rect 6884 -24770 6900 -24736
rect 7456 -24770 7472 -24736
rect 7902 -24770 7918 -24736
rect 8474 -24770 8490 -24736
rect 8920 -24770 8936 -24736
rect 9492 -24770 9508 -24736
rect 9938 -24770 9954 -24736
rect 10510 -24770 10526 -24736
rect 10956 -24770 10972 -24736
rect 11528 -24770 11544 -24736
rect 11974 -24770 11990 -24736
rect 12546 -24770 12562 -24736
rect 12992 -24770 13008 -24736
rect 13564 -24770 13580 -24736
rect 14010 -24770 14026 -24736
rect 14582 -24770 14598 -24736
rect 15028 -24770 15044 -24736
rect 15600 -24770 15616 -24736
rect 16046 -24770 16062 -24736
rect 16618 -24770 16634 -24736
rect 17064 -24770 17080 -24736
rect 17636 -24770 17652 -24736
rect 18082 -24770 18098 -24736
rect 18654 -24770 18670 -24736
rect 19100 -24770 19116 -24736
rect 19672 -24770 19688 -24736
rect 20118 -24770 20134 -24736
rect 20690 -24770 20706 -24736
rect 21136 -24770 21152 -24736
rect 21708 -24770 21724 -24736
rect 22154 -24770 22170 -24736
rect 22726 -24770 22742 -24736
rect -12322 -27222 -12222 -27060
rect 24822 -27222 24922 -27060
<< viali >>
rect 478 4222 540 4322
rect 540 4222 24660 4322
rect 24660 4222 24722 4322
rect 378 -9728 478 3702
rect 24722 -9728 24822 3702
rect 478 -10348 540 -10248
rect 540 -10348 24660 -10248
rect 24660 -10348 24722 -10248
rect -12222 -11278 -12160 -11178
rect -12160 -11278 24760 -11178
rect 24760 -11278 24822 -11178
rect -12322 -26330 -12222 -12070
rect -8890 -12474 -8426 -12440
rect -7872 -12474 -7408 -12440
rect -6854 -12474 -6390 -12440
rect -5836 -12474 -5372 -12440
rect -4818 -12474 -4354 -12440
rect -3800 -12474 -3336 -12440
rect -2782 -12474 -2318 -12440
rect -1764 -12474 -1300 -12440
rect -746 -12474 -282 -12440
rect -9184 -13100 -9150 -12524
rect -8166 -13100 -8132 -12524
rect -7148 -13100 -7114 -12524
rect -6130 -13100 -6096 -12524
rect -5112 -13100 -5078 -12524
rect -4094 -13100 -4060 -12524
rect -3076 -13100 -3042 -12524
rect -2058 -13100 -2024 -12524
rect -1040 -13100 -1006 -12524
rect -22 -13100 12 -12524
rect -8890 -13184 -8426 -13150
rect -7872 -13184 -7408 -13150
rect -6854 -13184 -6390 -13150
rect -5836 -13184 -5372 -13150
rect -4818 -13184 -4354 -13150
rect -3800 -13184 -3336 -13150
rect -2782 -13184 -2318 -13150
rect -1764 -13184 -1300 -13150
rect -746 -13184 -282 -13150
rect -8890 -13292 -8426 -13258
rect -7872 -13292 -7408 -13258
rect -6854 -13292 -6390 -13258
rect -5836 -13292 -5372 -13258
rect -4818 -13292 -4354 -13258
rect -3800 -13292 -3336 -13258
rect -2782 -13292 -2318 -13258
rect -1764 -13292 -1300 -13258
rect -746 -13292 -282 -13258
rect -9184 -13918 -9150 -13342
rect -8166 -13918 -8132 -13342
rect -7148 -13918 -7114 -13342
rect -6130 -13918 -6096 -13342
rect -5112 -13918 -5078 -13342
rect -4094 -13918 -4060 -13342
rect -3076 -13918 -3042 -13342
rect -2058 -13918 -2024 -13342
rect -1040 -13918 -1006 -13342
rect -22 -13918 12 -13342
rect -8890 -14002 -8426 -13968
rect -7872 -14002 -7408 -13968
rect -6854 -14002 -6390 -13968
rect -5836 -14002 -5372 -13968
rect -4818 -14002 -4354 -13968
rect -3800 -14002 -3336 -13968
rect -2782 -14002 -2318 -13968
rect -1764 -14002 -1300 -13968
rect -746 -14002 -282 -13968
rect -8890 -14110 -8426 -14076
rect -7872 -14110 -7408 -14076
rect -6854 -14110 -6390 -14076
rect -5836 -14110 -5372 -14076
rect -4818 -14110 -4354 -14076
rect -3800 -14110 -3336 -14076
rect -2782 -14110 -2318 -14076
rect -1764 -14110 -1300 -14076
rect -746 -14110 -282 -14076
rect -9184 -14736 -9150 -14160
rect -8166 -14736 -8132 -14160
rect -7148 -14736 -7114 -14160
rect -6130 -14736 -6096 -14160
rect -5112 -14736 -5078 -14160
rect -4094 -14736 -4060 -14160
rect -3076 -14736 -3042 -14160
rect -2058 -14736 -2024 -14160
rect -1040 -14736 -1006 -14160
rect -22 -14736 12 -14160
rect 2876 -14194 3340 -14160
rect 3894 -14194 4358 -14160
rect 4912 -14194 5376 -14160
rect 5930 -14194 6394 -14160
rect 6948 -14194 7412 -14160
rect 7966 -14194 8430 -14160
rect 8984 -14194 9448 -14160
rect 10002 -14194 10466 -14160
rect 11020 -14194 11484 -14160
rect 12038 -14194 12502 -14160
rect 13056 -14194 13520 -14160
rect 14074 -14194 14538 -14160
rect 15092 -14194 15556 -14160
rect 16110 -14194 16574 -14160
rect 17128 -14194 17592 -14160
rect 18146 -14194 18610 -14160
rect 19164 -14194 19628 -14160
rect 20182 -14194 20646 -14160
rect 21200 -14194 21664 -14160
rect 22218 -14194 22682 -14160
rect -8890 -14820 -8426 -14786
rect -7872 -14820 -7408 -14786
rect -6854 -14820 -6390 -14786
rect -5836 -14820 -5372 -14786
rect -4818 -14820 -4354 -14786
rect -3800 -14820 -3336 -14786
rect -2782 -14820 -2318 -14786
rect -1764 -14820 -1300 -14786
rect -746 -14820 -282 -14786
rect 2582 -14820 2616 -14244
rect 3600 -14820 3634 -14244
rect 4618 -14820 4652 -14244
rect 5636 -14820 5670 -14244
rect 6654 -14820 6688 -14244
rect 7672 -14820 7706 -14244
rect 8690 -14820 8724 -14244
rect 9708 -14820 9742 -14244
rect 10726 -14820 10760 -14244
rect 11744 -14820 11778 -14244
rect 12762 -14820 12796 -14244
rect 13780 -14820 13814 -14244
rect 14798 -14820 14832 -14244
rect 15816 -14820 15850 -14244
rect 16834 -14820 16868 -14244
rect 17852 -14820 17886 -14244
rect 18870 -14820 18904 -14244
rect 19888 -14820 19922 -14244
rect 20906 -14820 20940 -14244
rect 21924 -14820 21958 -14244
rect 22942 -14820 22976 -14244
rect -8890 -14928 -8426 -14894
rect -7872 -14928 -7408 -14894
rect -6854 -14928 -6390 -14894
rect -5836 -14928 -5372 -14894
rect -4818 -14928 -4354 -14894
rect -3800 -14928 -3336 -14894
rect -2782 -14928 -2318 -14894
rect -1764 -14928 -1300 -14894
rect -746 -14928 -282 -14894
rect 2876 -14904 3340 -14870
rect 3894 -14904 4358 -14870
rect 4912 -14904 5376 -14870
rect 5930 -14904 6394 -14870
rect 6948 -14904 7412 -14870
rect 7966 -14904 8430 -14870
rect 8984 -14904 9448 -14870
rect 10002 -14904 10466 -14870
rect 11020 -14904 11484 -14870
rect 12038 -14904 12502 -14870
rect 13056 -14904 13520 -14870
rect 14074 -14904 14538 -14870
rect 15092 -14904 15556 -14870
rect 16110 -14904 16574 -14870
rect 17128 -14904 17592 -14870
rect 18146 -14904 18610 -14870
rect 19164 -14904 19628 -14870
rect 20182 -14904 20646 -14870
rect 21200 -14904 21664 -14870
rect 22218 -14904 22682 -14870
rect -9184 -15554 -9150 -14978
rect -8166 -15554 -8132 -14978
rect -7148 -15554 -7114 -14978
rect -6130 -15554 -6096 -14978
rect -5112 -15554 -5078 -14978
rect -4094 -15554 -4060 -14978
rect -3076 -15554 -3042 -14978
rect -2058 -15554 -2024 -14978
rect -1040 -15554 -1006 -14978
rect -22 -15554 12 -14978
rect 2876 -15426 3340 -15392
rect 3894 -15426 4358 -15392
rect 4912 -15426 5376 -15392
rect 5930 -15426 6394 -15392
rect 6948 -15426 7412 -15392
rect 7966 -15426 8430 -15392
rect 8984 -15426 9448 -15392
rect 10002 -15426 10466 -15392
rect 11020 -15426 11484 -15392
rect 12038 -15426 12502 -15392
rect 13056 -15426 13520 -15392
rect 14074 -15426 14538 -15392
rect 15092 -15426 15556 -15392
rect 16110 -15426 16574 -15392
rect 17128 -15426 17592 -15392
rect 18146 -15426 18610 -15392
rect 19164 -15426 19628 -15392
rect 20182 -15426 20646 -15392
rect 21200 -15426 21664 -15392
rect 22218 -15426 22682 -15392
rect -8890 -15638 -8426 -15604
rect -7872 -15638 -7408 -15604
rect -6854 -15638 -6390 -15604
rect -5836 -15638 -5372 -15604
rect -4818 -15638 -4354 -15604
rect -3800 -15638 -3336 -15604
rect -2782 -15638 -2318 -15604
rect -1764 -15638 -1300 -15604
rect -746 -15638 -282 -15604
rect -8890 -15746 -8426 -15712
rect -7872 -15746 -7408 -15712
rect -6854 -15746 -6390 -15712
rect -5836 -15746 -5372 -15712
rect -4818 -15746 -4354 -15712
rect -3800 -15746 -3336 -15712
rect -2782 -15746 -2318 -15712
rect -1764 -15746 -1300 -15712
rect -746 -15746 -282 -15712
rect -9184 -16372 -9150 -15796
rect -8166 -16372 -8132 -15796
rect -7148 -16372 -7114 -15796
rect -6130 -16372 -6096 -15796
rect -5112 -16372 -5078 -15796
rect -4094 -16372 -4060 -15796
rect -3076 -16372 -3042 -15796
rect -2058 -16372 -2024 -15796
rect -1040 -16372 -1006 -15796
rect -22 -16372 12 -15796
rect 2582 -16052 2616 -15476
rect 3600 -16052 3634 -15476
rect 4618 -16052 4652 -15476
rect 5636 -16052 5670 -15476
rect 6654 -16052 6688 -15476
rect 7672 -16052 7706 -15476
rect 8690 -16052 8724 -15476
rect 9708 -16052 9742 -15476
rect 10726 -16052 10760 -15476
rect 11744 -16052 11778 -15476
rect 12762 -16052 12796 -15476
rect 13780 -16052 13814 -15476
rect 14798 -16052 14832 -15476
rect 15816 -16052 15850 -15476
rect 16834 -16052 16868 -15476
rect 17852 -16052 17886 -15476
rect 18870 -16052 18904 -15476
rect 19888 -16052 19922 -15476
rect 20906 -16052 20940 -15476
rect 21924 -16052 21958 -15476
rect 22942 -16052 22976 -15476
rect 2876 -16136 3340 -16102
rect 3894 -16136 4358 -16102
rect 4912 -16136 5376 -16102
rect 5930 -16136 6394 -16102
rect 6948 -16136 7412 -16102
rect 7966 -16136 8430 -16102
rect 8984 -16136 9448 -16102
rect 10002 -16136 10466 -16102
rect 11020 -16136 11484 -16102
rect 12038 -16136 12502 -16102
rect 13056 -16136 13520 -16102
rect 14074 -16136 14538 -16102
rect 15092 -16136 15556 -16102
rect 16110 -16136 16574 -16102
rect 17128 -16134 17592 -16102
rect 17128 -16136 17318 -16134
rect 17378 -16136 17592 -16134
rect 18146 -16130 18610 -16102
rect 18146 -16136 18352 -16130
rect 18412 -16136 18610 -16130
rect 19164 -16136 19628 -16102
rect 20182 -16136 20646 -16102
rect 21200 -16136 21664 -16102
rect 22218 -16136 22682 -16102
rect -8890 -16456 -8426 -16422
rect -7872 -16456 -7408 -16422
rect -6854 -16456 -6390 -16422
rect -5836 -16456 -5372 -16422
rect -4818 -16456 -4354 -16422
rect -3800 -16456 -3336 -16422
rect -2782 -16456 -2318 -16422
rect -1764 -16456 -1300 -16422
rect -746 -16456 -282 -16422
rect -8890 -16564 -8426 -16530
rect -7872 -16564 -7408 -16530
rect -6854 -16564 -6390 -16530
rect -5836 -16564 -5372 -16530
rect -4818 -16564 -4354 -16530
rect -3800 -16564 -3336 -16530
rect -2782 -16564 -2318 -16530
rect -1764 -16564 -1300 -16530
rect -746 -16564 -282 -16530
rect -9184 -17190 -9150 -16614
rect -8166 -17190 -8132 -16614
rect -7148 -17190 -7114 -16614
rect -6130 -17190 -6096 -16614
rect -5112 -17190 -5078 -16614
rect -4094 -17190 -4060 -16614
rect -3076 -17190 -3042 -16614
rect -2058 -17190 -2024 -16614
rect -1040 -17190 -1006 -16614
rect -22 -17190 12 -16614
rect 2874 -16660 3338 -16626
rect 3892 -16660 4356 -16626
rect 4910 -16660 5374 -16626
rect 5928 -16660 6392 -16626
rect 6946 -16660 7410 -16626
rect 7964 -16660 8428 -16626
rect 8982 -16660 9446 -16626
rect 10000 -16660 10464 -16626
rect 11018 -16660 11482 -16626
rect 12036 -16660 12500 -16626
rect 13054 -16660 13518 -16626
rect 14072 -16660 14536 -16626
rect 15090 -16660 15554 -16626
rect 16108 -16660 16572 -16626
rect 17126 -16660 17590 -16626
rect 18144 -16660 18608 -16626
rect 19162 -16660 19626 -16626
rect 20180 -16660 20644 -16626
rect 21198 -16660 21662 -16626
rect 22216 -16660 22680 -16626
rect -8890 -17274 -8426 -17240
rect -7872 -17274 -7408 -17240
rect -6854 -17274 -6390 -17240
rect -5836 -17274 -5372 -17240
rect -4818 -17274 -4354 -17240
rect -3800 -17274 -3336 -17240
rect -2782 -17274 -2318 -17240
rect -1764 -17274 -1300 -17240
rect -746 -17274 -282 -17240
rect 2580 -17286 2614 -16710
rect 3598 -17286 3632 -16710
rect 4616 -17286 4650 -16710
rect 5634 -17286 5668 -16710
rect 6652 -17286 6686 -16710
rect 7670 -17286 7704 -16710
rect 8688 -17286 8722 -16710
rect 9706 -17286 9740 -16710
rect 10724 -17286 10758 -16710
rect 11742 -17286 11776 -16710
rect 12760 -17286 12794 -16710
rect 13778 -17286 13812 -16710
rect 14796 -17286 14830 -16710
rect 15814 -17286 15848 -16710
rect 16832 -17286 16866 -16710
rect 17850 -17286 17884 -16710
rect 18868 -17286 18902 -16710
rect 19886 -17286 19920 -16710
rect 20904 -17286 20938 -16710
rect 21922 -17286 21956 -16710
rect 22940 -17286 22974 -16710
rect -8890 -17382 -8426 -17348
rect -7872 -17382 -7408 -17348
rect -6854 -17382 -6390 -17348
rect -5836 -17382 -5372 -17348
rect -4818 -17382 -4354 -17348
rect -3800 -17382 -3336 -17348
rect -2782 -17382 -2318 -17348
rect -1764 -17382 -1300 -17348
rect -746 -17382 -282 -17348
rect 2874 -17370 3338 -17336
rect 3892 -17370 4356 -17336
rect 4910 -17370 5374 -17336
rect 5928 -17370 6392 -17336
rect 6946 -17370 7410 -17336
rect 7964 -17370 8428 -17336
rect 8982 -17370 9446 -17336
rect 10000 -17370 10464 -17336
rect 11018 -17370 11482 -17336
rect 12036 -17370 12500 -17336
rect 13054 -17370 13518 -17336
rect 14072 -17370 14536 -17336
rect 15090 -17370 15554 -17336
rect 16108 -17370 16572 -17336
rect 17126 -17370 17590 -17336
rect 18144 -17370 18608 -17336
rect 19162 -17370 19626 -17336
rect 20180 -17370 20644 -17336
rect 21198 -17370 21662 -17336
rect 22216 -17370 22680 -17336
rect -9184 -18008 -9150 -17432
rect -8166 -18008 -8132 -17432
rect -7148 -18008 -7114 -17432
rect -6130 -18008 -6096 -17432
rect -5112 -18008 -5078 -17432
rect -4094 -18008 -4060 -17432
rect -3076 -18008 -3042 -17432
rect -2058 -18008 -2024 -17432
rect -1040 -18008 -1006 -17432
rect -22 -18008 12 -17432
rect 2874 -17894 3338 -17860
rect 3892 -17894 4356 -17860
rect 4910 -17894 5374 -17860
rect 5928 -17894 6392 -17860
rect 6946 -17894 7410 -17860
rect 7964 -17894 8428 -17860
rect 8982 -17894 9446 -17860
rect 10000 -17894 10464 -17860
rect 11018 -17894 11482 -17860
rect 12036 -17894 12500 -17860
rect 13054 -17894 13518 -17860
rect 14072 -17894 14536 -17860
rect 15090 -17894 15554 -17860
rect 16108 -17894 16572 -17860
rect 17126 -17894 17590 -17860
rect 18144 -17894 18608 -17860
rect 19162 -17894 19626 -17860
rect 20180 -17894 20644 -17860
rect 21198 -17894 21662 -17860
rect 22216 -17894 22680 -17860
rect -8890 -18092 -8426 -18058
rect -7872 -18092 -7408 -18058
rect -6854 -18092 -6390 -18058
rect -5836 -18092 -5372 -18058
rect -4818 -18092 -4354 -18058
rect -3800 -18092 -3336 -18058
rect -2782 -18092 -2318 -18058
rect -1764 -18092 -1300 -18058
rect -746 -18092 -282 -18058
rect -8890 -18200 -8426 -18166
rect -7872 -18200 -7408 -18166
rect -6854 -18200 -6390 -18166
rect -5836 -18200 -5372 -18166
rect -4818 -18200 -4354 -18166
rect -3800 -18200 -3336 -18166
rect -2782 -18200 -2318 -18166
rect -1764 -18200 -1300 -18166
rect -746 -18200 -282 -18166
rect -9184 -18826 -9150 -18250
rect -8166 -18826 -8132 -18250
rect -7148 -18826 -7114 -18250
rect -6130 -18826 -6096 -18250
rect -5112 -18826 -5078 -18250
rect -4094 -18826 -4060 -18250
rect -3076 -18826 -3042 -18250
rect -2058 -18826 -2024 -18250
rect -1040 -18826 -1006 -18250
rect -22 -18826 12 -18250
rect 2580 -18520 2614 -17944
rect 3598 -18520 3632 -17944
rect 4616 -18520 4650 -17944
rect 5634 -18520 5668 -17944
rect 6652 -18520 6686 -17944
rect 7670 -18520 7704 -17944
rect 8688 -18520 8722 -17944
rect 9706 -18520 9740 -17944
rect 10724 -18520 10758 -17944
rect 11742 -18520 11776 -17944
rect 12760 -18520 12794 -17944
rect 13778 -18520 13812 -17944
rect 14796 -18520 14830 -17944
rect 15814 -18520 15848 -17944
rect 16832 -18520 16866 -17944
rect 17850 -18520 17884 -17944
rect 18868 -18520 18902 -17944
rect 19886 -18520 19920 -17944
rect 20904 -18520 20938 -17944
rect 21922 -18520 21956 -17944
rect 22940 -18520 22974 -17944
rect 2874 -18604 3338 -18570
rect 3892 -18604 4356 -18570
rect 4910 -18604 5374 -18570
rect 5928 -18604 6392 -18570
rect 6946 -18604 7410 -18570
rect 7964 -18604 8428 -18570
rect 8982 -18604 9446 -18570
rect 10000 -18604 10464 -18570
rect 11018 -18604 11482 -18570
rect 12036 -18604 12500 -18570
rect 13054 -18604 13518 -18570
rect 14072 -18604 14536 -18570
rect 15090 -18604 15554 -18570
rect 16108 -18604 16572 -18570
rect 17126 -18604 17590 -18570
rect 18144 -18604 18608 -18570
rect 19162 -18604 19626 -18570
rect 20180 -18604 20644 -18570
rect 21198 -18604 21662 -18570
rect 22216 -18604 22680 -18570
rect -8890 -18910 -8426 -18876
rect -7872 -18910 -7408 -18876
rect -6854 -18910 -6390 -18876
rect -5836 -18910 -5372 -18876
rect -4818 -18910 -4354 -18876
rect -3800 -18910 -3336 -18876
rect -2782 -18910 -2318 -18876
rect -1764 -18910 -1300 -18876
rect -746 -18910 -282 -18876
rect 2874 -19126 3338 -19092
rect 3892 -19126 4356 -19092
rect 4910 -19126 5374 -19092
rect 5928 -19126 6392 -19092
rect 6946 -19126 7410 -19092
rect 7964 -19126 8428 -19092
rect 8982 -19126 9446 -19092
rect 10000 -19126 10464 -19092
rect 11018 -19126 11482 -19092
rect 12036 -19126 12500 -19092
rect 13054 -19126 13518 -19092
rect 14072 -19126 14536 -19092
rect 15090 -19126 15554 -19092
rect 16108 -19126 16572 -19092
rect 17126 -19126 17590 -19092
rect 18144 -19126 18608 -19092
rect 19162 -19126 19626 -19092
rect 20180 -19126 20644 -19092
rect 21198 -19126 21662 -19092
rect 22216 -19126 22680 -19092
rect 2580 -19752 2614 -19176
rect 3598 -19752 3632 -19176
rect 4616 -19752 4650 -19176
rect 5634 -19752 5668 -19176
rect 6652 -19752 6686 -19176
rect 7670 -19752 7704 -19176
rect 8688 -19752 8722 -19176
rect 9706 -19752 9740 -19176
rect 10724 -19752 10758 -19176
rect 11742 -19752 11776 -19176
rect 12760 -19752 12794 -19176
rect 13778 -19752 13812 -19176
rect 14796 -19752 14830 -19176
rect 15814 -19752 15848 -19176
rect 16832 -19752 16866 -19176
rect 17850 -19752 17884 -19176
rect 18868 -19752 18902 -19176
rect 19886 -19752 19920 -19176
rect 20904 -19752 20938 -19176
rect 21922 -19752 21956 -19176
rect 22940 -19752 22974 -19176
rect 2874 -19836 3338 -19802
rect 3892 -19836 4356 -19802
rect 4910 -19836 5374 -19802
rect 5928 -19836 6392 -19802
rect 6946 -19836 7410 -19802
rect 7964 -19836 8428 -19802
rect 8982 -19836 9446 -19802
rect 10000 -19836 10464 -19802
rect 11018 -19836 11482 -19802
rect 12036 -19836 12500 -19802
rect 13054 -19836 13518 -19802
rect 14072 -19836 14536 -19802
rect 15090 -19836 15554 -19802
rect 16108 -19836 16572 -19802
rect 17126 -19836 17590 -19802
rect 18144 -19836 18608 -19802
rect 19162 -19836 19626 -19802
rect 20180 -19836 20644 -19802
rect 21198 -19836 21662 -19802
rect 22216 -19836 22680 -19802
rect 2874 -20360 3338 -20326
rect 3892 -20360 4356 -20326
rect 4910 -20360 5374 -20326
rect 5928 -20360 6392 -20326
rect 6946 -20360 7410 -20326
rect 7964 -20360 8428 -20326
rect 8982 -20360 9446 -20326
rect 10000 -20360 10464 -20326
rect 11018 -20360 11482 -20326
rect 12036 -20360 12500 -20326
rect 13054 -20360 13518 -20326
rect 14072 -20360 14536 -20326
rect 15090 -20360 15554 -20326
rect 16108 -20360 16572 -20326
rect 17126 -20360 17590 -20326
rect 18144 -20360 18608 -20326
rect 19162 -20360 19626 -20326
rect 20180 -20360 20644 -20326
rect 21198 -20360 21662 -20326
rect 22216 -20360 22680 -20326
rect 2580 -20986 2614 -20410
rect 3598 -20986 3632 -20410
rect 4616 -20986 4650 -20410
rect 5634 -20986 5668 -20410
rect 6652 -20986 6686 -20410
rect 7670 -20986 7704 -20410
rect 8688 -20986 8722 -20410
rect 9706 -20986 9740 -20410
rect 10724 -20986 10758 -20410
rect 11742 -20986 11776 -20410
rect 12760 -20986 12794 -20410
rect 13778 -20986 13812 -20410
rect 14796 -20986 14830 -20410
rect 15814 -20986 15848 -20410
rect 16832 -20986 16866 -20410
rect 17850 -20986 17884 -20410
rect 18868 -20986 18902 -20410
rect 19886 -20986 19920 -20410
rect 20904 -20986 20938 -20410
rect 21922 -20986 21956 -20410
rect 22940 -20986 22974 -20410
rect 2874 -21070 3338 -21036
rect 3892 -21070 4356 -21036
rect 4910 -21070 5374 -21036
rect 5928 -21070 6392 -21036
rect 6946 -21070 7410 -21036
rect 7964 -21070 8428 -21036
rect 8982 -21070 9446 -21036
rect 10000 -21070 10464 -21036
rect 11018 -21070 11482 -21036
rect 12036 -21070 12500 -21036
rect 13054 -21070 13518 -21036
rect 14072 -21070 14536 -21036
rect 15090 -21070 15554 -21036
rect 16108 -21070 16572 -21036
rect 17126 -21070 17590 -21036
rect 18144 -21070 18608 -21036
rect 19162 -21070 19626 -21036
rect 20180 -21070 20644 -21036
rect 21198 -21070 21662 -21036
rect 22216 -21070 22680 -21036
rect 2874 -21594 3338 -21560
rect 3892 -21594 4356 -21560
rect 4910 -21594 5374 -21560
rect 5928 -21594 6392 -21560
rect 6946 -21594 7410 -21560
rect 7964 -21594 8428 -21560
rect 8982 -21594 9446 -21560
rect 10000 -21594 10464 -21560
rect 11018 -21594 11482 -21560
rect 12036 -21594 12500 -21560
rect 13054 -21594 13518 -21560
rect 14072 -21594 14536 -21560
rect 15090 -21594 15554 -21560
rect 16108 -21594 16572 -21560
rect 17126 -21594 17590 -21560
rect 18144 -21594 18608 -21560
rect 19162 -21594 19626 -21560
rect 20180 -21594 20644 -21560
rect 21198 -21594 21662 -21560
rect 22216 -21594 22680 -21560
rect 2580 -22220 2614 -21644
rect 3598 -22220 3632 -21644
rect 4616 -22220 4650 -21644
rect 5634 -22220 5668 -21644
rect 6652 -22220 6686 -21644
rect 7670 -22220 7704 -21644
rect 8688 -22220 8722 -21644
rect 9706 -22220 9740 -21644
rect 10724 -22220 10758 -21644
rect 11742 -22220 11776 -21644
rect 12760 -22220 12794 -21644
rect 13778 -22220 13812 -21644
rect 14796 -22220 14830 -21644
rect 15814 -22220 15848 -21644
rect 16832 -22220 16866 -21644
rect 17850 -22220 17884 -21644
rect 18868 -22220 18902 -21644
rect 19886 -22220 19920 -21644
rect 20904 -22220 20938 -21644
rect 21922 -22220 21956 -21644
rect 22940 -22220 22974 -21644
rect 2874 -22304 3338 -22270
rect 3892 -22304 4356 -22270
rect 4910 -22304 5374 -22270
rect 5928 -22304 6392 -22270
rect 6946 -22304 7410 -22270
rect 7964 -22304 8428 -22270
rect 8982 -22304 9446 -22270
rect 10000 -22304 10464 -22270
rect 11018 -22304 11482 -22270
rect 12036 -22304 12500 -22270
rect 13054 -22304 13518 -22270
rect 14072 -22304 14536 -22270
rect 15090 -22304 15554 -22270
rect 16108 -22304 16572 -22270
rect 17126 -22304 17590 -22270
rect 18144 -22304 18608 -22270
rect 19162 -22304 19626 -22270
rect 20180 -22304 20644 -22270
rect 21198 -22304 21662 -22270
rect 22216 -22304 22680 -22270
rect 2874 -22826 3338 -22792
rect 3892 -22826 4356 -22792
rect 4910 -22826 5374 -22792
rect 5928 -22826 6392 -22792
rect 6946 -22826 7410 -22792
rect 7964 -22826 8428 -22792
rect 8982 -22826 9446 -22792
rect 10000 -22826 10464 -22792
rect 11018 -22826 11482 -22792
rect 12036 -22826 12500 -22792
rect 13054 -22826 13518 -22792
rect 14072 -22826 14536 -22792
rect 15090 -22826 15554 -22792
rect 16108 -22826 16572 -22792
rect 17126 -22826 17590 -22792
rect 18144 -22826 18608 -22792
rect 19162 -22826 19626 -22792
rect 20180 -22826 20644 -22792
rect 21198 -22826 21662 -22792
rect 22216 -22826 22680 -22792
rect 2580 -23452 2614 -22876
rect 3598 -23452 3632 -22876
rect 4616 -23452 4650 -22876
rect 5634 -23452 5668 -22876
rect 6652 -23452 6686 -22876
rect 7670 -23452 7704 -22876
rect 8688 -23452 8722 -22876
rect 9706 -23452 9740 -22876
rect 10724 -23452 10758 -22876
rect 11742 -23452 11776 -22876
rect 12760 -23452 12794 -22876
rect 13778 -23452 13812 -22876
rect 14796 -23452 14830 -22876
rect 15814 -23452 15848 -22876
rect 16832 -23452 16866 -22876
rect 17850 -23452 17884 -22876
rect 18868 -23452 18902 -22876
rect 19886 -23452 19920 -22876
rect 20904 -23452 20938 -22876
rect 21922 -23452 21956 -22876
rect 22940 -23452 22974 -22876
rect 2874 -23536 3338 -23502
rect 3892 -23536 4356 -23502
rect 4910 -23536 5374 -23502
rect 5928 -23536 6392 -23502
rect 6946 -23536 7410 -23502
rect 7964 -23536 8428 -23502
rect 8982 -23536 9446 -23502
rect 10000 -23536 10464 -23502
rect 11018 -23536 11482 -23502
rect 12036 -23536 12500 -23502
rect 13054 -23536 13518 -23502
rect 14072 -23536 14536 -23502
rect 15090 -23536 15554 -23502
rect 16108 -23536 16572 -23502
rect 17126 -23536 17590 -23502
rect 18144 -23536 18608 -23502
rect 19162 -23536 19626 -23502
rect 20180 -23536 20644 -23502
rect 21198 -23536 21662 -23502
rect 22216 -23536 22680 -23502
rect 2874 -24060 3338 -24026
rect 3892 -24060 4356 -24026
rect 4910 -24060 5374 -24026
rect 5928 -24060 6392 -24026
rect 6946 -24060 7410 -24026
rect 7964 -24060 8428 -24026
rect 8982 -24060 9446 -24026
rect 10000 -24060 10464 -24026
rect 11018 -24060 11482 -24026
rect 12036 -24060 12500 -24026
rect 13054 -24060 13518 -24026
rect 14072 -24060 14536 -24026
rect 15090 -24060 15554 -24026
rect 16108 -24060 16572 -24026
rect 17126 -24060 17590 -24026
rect 18144 -24060 18608 -24026
rect 19162 -24060 19626 -24026
rect 20180 -24060 20644 -24026
rect 21198 -24060 21662 -24026
rect 22216 -24060 22680 -24026
rect 2580 -24686 2614 -24110
rect 3598 -24686 3632 -24110
rect 4616 -24686 4650 -24110
rect 5634 -24686 5668 -24110
rect 6652 -24686 6686 -24110
rect 7670 -24686 7704 -24110
rect 8688 -24686 8722 -24110
rect 9706 -24686 9740 -24110
rect 10724 -24686 10758 -24110
rect 11742 -24686 11776 -24110
rect 12760 -24686 12794 -24110
rect 13778 -24686 13812 -24110
rect 14796 -24686 14830 -24110
rect 15814 -24686 15848 -24110
rect 16832 -24686 16866 -24110
rect 17850 -24686 17884 -24110
rect 18868 -24686 18902 -24110
rect 19886 -24686 19920 -24110
rect 20904 -24686 20938 -24110
rect 21922 -24686 21956 -24110
rect 22940 -24686 22974 -24110
rect 2874 -24770 3338 -24736
rect 3892 -24770 4356 -24736
rect 4910 -24770 5374 -24736
rect 5928 -24770 6392 -24736
rect 6946 -24770 7410 -24736
rect 7964 -24770 8428 -24736
rect 8982 -24770 9446 -24736
rect 10000 -24770 10464 -24736
rect 11018 -24770 11482 -24736
rect 12036 -24770 12500 -24736
rect 13054 -24770 13518 -24736
rect 14072 -24770 14536 -24736
rect 15090 -24770 15554 -24736
rect 16108 -24770 16572 -24736
rect 17126 -24770 17590 -24736
rect 18144 -24770 18608 -24736
rect 19162 -24770 19626 -24736
rect 20180 -24770 20644 -24736
rect 21198 -24770 21662 -24736
rect 22216 -24770 22680 -24736
rect 24822 -26330 24922 -12070
rect -12222 -27222 -12160 -27122
rect -12160 -27222 24760 -27122
rect 24760 -27222 24822 -27122
<< metal1 >>
rect 372 4322 24828 4328
rect 372 4222 478 4322
rect 24722 4222 24828 4322
rect 372 4216 24828 4222
rect 372 3702 484 4216
rect 1084 3916 1094 4216
rect 24106 3916 24116 4216
rect 372 -9728 378 3702
rect 478 -9728 484 3702
rect 3998 3834 20878 3866
rect 3998 3620 4061 3834
rect 20846 3620 20878 3834
rect 3998 3598 4048 3620
rect 4108 3598 4484 3620
rect 4544 3598 4922 3620
rect 4982 3598 5356 3620
rect 5416 3600 20878 3620
rect 24716 3702 24828 4216
rect 5416 3598 8352 3600
rect 8512 2124 8572 3600
rect 10548 2124 10608 3600
rect 11052 2124 11112 3600
rect 11560 2124 11620 3600
rect 12072 2124 12132 3600
rect 12586 2124 12646 3600
rect 14618 2124 14678 3600
rect 16658 2124 16718 3600
rect 17148 2124 17208 3600
rect 17668 2124 17728 3600
rect 18176 2124 18236 3600
rect 18690 2124 18750 3600
rect 20726 2124 20786 3600
rect 8512 2064 20786 2124
rect 7980 1858 7986 1918
rect 8046 1858 8052 1918
rect 6474 1642 7552 1702
rect 6474 1422 6534 1642
rect 6978 1526 7038 1642
rect 7492 1436 7552 1642
rect 7986 1518 8046 1858
rect 8512 1672 8572 2064
rect 9062 1858 9068 1918
rect 9128 1858 9134 1918
rect 10020 1858 10026 1918
rect 10086 1858 10092 1918
rect 8506 1612 8512 1672
rect 8572 1612 8578 1672
rect 8512 1438 8572 1612
rect 9068 1516 9128 1858
rect 10026 1512 10086 1858
rect 10548 1672 10608 2064
rect 10542 1612 10548 1672
rect 10608 1612 10614 1672
rect 10548 1438 10608 1612
rect 11052 1518 11112 2064
rect 11560 1392 11620 2064
rect 12072 1518 12132 2064
rect 12586 1674 12646 2064
rect 13084 1858 13090 1918
rect 13150 1858 13156 1918
rect 14102 1858 14108 1918
rect 14168 1858 14174 1918
rect 12580 1614 12586 1674
rect 12646 1614 12652 1674
rect 12586 1422 12646 1614
rect 13090 1522 13150 1858
rect 14108 1516 14168 1858
rect 14618 1674 14678 2064
rect 15126 1858 15132 1918
rect 15192 1858 15198 1918
rect 16138 1858 16144 1918
rect 16204 1858 16210 1918
rect 14610 1614 14616 1674
rect 14676 1614 14682 1674
rect 14618 1422 14678 1614
rect 15132 1522 15192 1858
rect 16144 1522 16204 1858
rect 16658 1676 16718 2064
rect 16652 1616 16658 1676
rect 16718 1616 16724 1676
rect 16658 1424 16718 1616
rect 17148 1522 17208 2064
rect 17668 1676 17728 2064
rect 17662 1616 17668 1676
rect 17728 1616 17734 1676
rect 17668 1392 17728 1616
rect 18176 1512 18236 2064
rect 18690 1676 18750 2064
rect 19196 1858 19202 1918
rect 19262 1858 19268 1918
rect 20208 1858 20214 1918
rect 20274 1858 20280 1918
rect 18684 1616 18690 1676
rect 18750 1616 18756 1676
rect 18690 1434 18750 1616
rect 19202 1522 19262 1858
rect 20214 1522 20274 1858
rect 20726 1676 20786 2064
rect 21226 1858 21232 1918
rect 21292 1858 21298 1918
rect 20720 1616 20726 1676
rect 20786 1616 20792 1676
rect 20726 1430 20786 1616
rect 21232 1516 21292 1858
rect 21746 1624 22826 1684
rect 21746 1432 21806 1624
rect 22248 1522 22308 1624
rect 22766 1416 22826 1624
rect 7494 740 7554 922
rect 6324 680 6330 740
rect 6390 680 6396 740
rect 7488 680 7494 740
rect 7554 680 7560 740
rect 6194 476 6200 536
rect 6260 476 6266 536
rect 4186 -1708 4192 -1648
rect 4252 -1708 4258 -1648
rect 2014 -5024 3236 -4964
rect 2014 -6940 2074 -5024
rect 2156 -5238 2216 -5024
rect 2668 -5128 2728 -5024
rect 3176 -5240 3236 -5024
rect 3676 -5906 3736 -5824
rect 3670 -5966 3676 -5906
rect 3736 -5966 3742 -5906
rect 3778 -6078 3784 -6018
rect 3844 -6078 3850 -6018
rect 3784 -6158 3844 -6078
rect 2008 -7000 2014 -6940
rect 2074 -7000 2080 -6940
rect 1888 -8028 1948 -8022
rect 2014 -8028 2074 -7000
rect 2154 -7050 2214 -6738
rect 2656 -7050 2716 -6856
rect 3174 -7050 3234 -6746
rect 2154 -7110 3174 -7050
rect 3234 -7110 3240 -7050
rect 2154 -7312 2214 -7110
rect 2656 -7188 2716 -7110
rect 3174 -7316 3234 -7110
rect 3684 -7194 3744 -6860
rect 3690 -7974 3750 -7888
rect 1948 -8088 3238 -8028
rect 3684 -8034 3690 -7974
rect 3750 -8034 3756 -7974
rect 1888 -8094 1948 -8088
rect 2152 -8336 2212 -8088
rect 2660 -8226 2720 -8088
rect 3178 -8332 3238 -8088
rect 3790 -8134 3796 -8074
rect 3856 -8134 3862 -8074
rect 3796 -8222 3856 -8134
rect 4192 -8358 4252 -1708
rect 6200 -2080 6260 476
rect 6330 -1934 6390 680
rect 7488 476 7494 536
rect 7554 476 7560 536
rect 7494 288 7554 476
rect 7998 376 8058 834
rect 8514 286 8574 926
rect 9530 636 9590 914
rect 9524 576 9530 636
rect 9590 576 9596 636
rect 10538 296 10602 944
rect 11560 576 11566 636
rect 11626 576 11632 636
rect 11566 288 11626 576
rect 12574 292 12638 940
rect 13092 378 13152 836
rect 13604 740 13664 926
rect 13598 680 13604 740
rect 13664 680 13670 740
rect 13594 476 13600 536
rect 13660 476 13666 536
rect 13600 300 13660 476
rect 14110 384 14170 842
rect 14616 294 14680 942
rect 15126 376 15186 839
rect 15638 740 15698 924
rect 15632 680 15638 740
rect 15698 680 15704 740
rect 16138 536 16198 839
rect 15630 476 15636 536
rect 15696 476 15702 536
rect 16132 476 16138 536
rect 16198 476 16204 536
rect 15636 294 15696 476
rect 16138 376 16198 476
rect 16654 278 16718 926
rect 17666 576 17672 636
rect 17732 576 17738 636
rect 17152 476 17158 536
rect 17218 476 17224 536
rect 17158 382 17218 476
rect 17672 302 17732 576
rect 18178 476 18184 536
rect 18244 476 18250 536
rect 18690 532 18750 934
rect 19706 636 19766 918
rect 19700 576 19706 636
rect 19766 576 19772 636
rect 20730 538 20790 924
rect 20730 532 20794 538
rect 18184 382 18244 476
rect 18684 472 18690 532
rect 18750 472 18756 532
rect 19198 472 19204 532
rect 19264 472 19270 532
rect 19702 472 19708 532
rect 19768 472 19774 532
rect 20208 472 20214 532
rect 20274 472 20280 532
rect 20730 472 20734 532
rect 18690 282 18750 472
rect 19204 380 19264 472
rect 19708 298 19768 472
rect 20214 380 20274 472
rect 20730 466 20794 472
rect 20730 290 20790 466
rect 21210 382 21270 845
rect 21746 740 21806 926
rect 21740 680 21746 740
rect 21806 680 21812 740
rect 22990 680 22996 740
rect 23056 680 23062 740
rect 21750 464 22820 524
rect 21750 298 21810 464
rect 22256 390 22316 464
rect 22760 292 22820 464
rect 14618 -204 14678 -202
rect 6476 -400 6536 -214
rect 6988 -400 7048 -312
rect 7494 -400 7554 -220
rect 10546 -224 10606 -222
rect 6476 -460 7554 -400
rect 7488 -604 7548 -602
rect 6478 -664 7548 -604
rect 6478 -842 6538 -664
rect 6988 -744 7048 -664
rect 7488 -842 7548 -664
rect 7980 -614 8040 -296
rect 7980 -754 8040 -674
rect 8510 -396 8570 -224
rect 9008 -396 9068 -302
rect 9528 -396 9588 -230
rect 10036 -396 10096 -298
rect 8510 -398 10096 -396
rect 10546 -398 10610 -224
rect 8510 -456 10036 -398
rect 8510 -862 8570 -456
rect 10540 -458 10546 -398
rect 10606 -458 10612 -398
rect 10036 -464 10096 -458
rect 9522 -560 9528 -496
rect 9592 -560 9598 -496
rect 9012 -674 9018 -614
rect 9078 -674 9084 -614
rect 9528 -654 9592 -560
rect 9018 -754 9078 -674
rect 9528 -856 9594 -654
rect 10024 -674 10030 -614
rect 10090 -674 10096 -614
rect 10030 -758 10090 -674
rect 9528 -860 9592 -856
rect 10546 -858 10610 -458
rect 11040 -606 11100 -310
rect 11564 -496 11628 -214
rect 12580 -216 12640 -214
rect 11398 -560 11404 -496
rect 11468 -560 11628 -496
rect 12064 -606 12124 -310
rect 12580 -398 12644 -216
rect 12574 -458 12580 -398
rect 12640 -458 12646 -398
rect 11034 -666 11040 -606
rect 11100 -666 11106 -606
rect 12058 -666 12064 -606
rect 12124 -666 12130 -606
rect 12580 -870 12644 -458
rect 13092 -606 13152 -296
rect 13086 -666 13092 -606
rect 13152 -666 13158 -606
rect 13092 -754 13152 -666
rect 14120 -764 14180 -306
rect 14618 -400 14682 -204
rect 16654 -208 16714 -206
rect 14612 -460 14618 -400
rect 14678 -460 14684 -400
rect 14618 -850 14682 -460
rect 15138 -754 15198 -291
rect 15638 -498 15698 -220
rect 15632 -558 15638 -498
rect 15698 -558 15704 -498
rect 16138 -758 16198 -295
rect 16654 -400 16718 -208
rect 18690 -400 18750 -214
rect 19192 -400 19252 -308
rect 16648 -460 16654 -400
rect 16714 -460 16720 -400
rect 17148 -460 17154 -400
rect 17214 -460 17220 -400
rect 17662 -460 17668 -400
rect 17728 -460 17734 -400
rect 18186 -460 18192 -400
rect 18252 -460 18258 -400
rect 18684 -460 18690 -400
rect 18750 -460 18756 -400
rect 19186 -460 19192 -400
rect 19252 -460 19258 -400
rect 19706 -402 19766 -180
rect 20724 -220 20784 -218
rect 20214 -402 20274 -296
rect 20724 -402 20788 -220
rect 16654 -862 16718 -460
rect 17154 -754 17214 -460
rect 17668 -864 17728 -460
rect 18192 -754 18252 -460
rect 18690 -864 18750 -460
rect 19700 -462 19706 -402
rect 19766 -462 19772 -402
rect 20208 -462 20214 -402
rect 20274 -462 20280 -402
rect 20718 -462 20724 -402
rect 20784 -462 20790 -402
rect 19190 -674 19196 -614
rect 19256 -674 19262 -614
rect 20202 -674 20208 -614
rect 20268 -674 20274 -614
rect 19196 -756 19256 -674
rect 20208 -750 20268 -674
rect 20724 -856 20788 -462
rect 21210 -614 21270 -297
rect 21746 -498 21806 -220
rect 21740 -558 21746 -498
rect 21806 -558 21812 -498
rect 21748 -612 21808 -610
rect 21204 -674 21210 -614
rect 21270 -674 21276 -614
rect 21748 -672 22820 -612
rect 21210 -760 21270 -674
rect 21748 -836 21808 -672
rect 22252 -748 22312 -672
rect 22760 -860 22820 -672
rect 7488 -1594 7552 -1344
rect 7044 -1654 7552 -1594
rect 6324 -1994 6330 -1934
rect 6390 -1994 6396 -1934
rect 6200 -2140 6620 -2080
rect 6560 -4952 6620 -2140
rect 6680 -4402 6686 -4342
rect 6746 -4402 6752 -4342
rect 5210 -5020 6420 -4960
rect 6554 -5012 6560 -4952
rect 6620 -5012 6626 -4952
rect 5210 -5236 5270 -5020
rect 5722 -5124 5782 -5020
rect 6228 -5234 6288 -5020
rect 4568 -6018 4628 -5822
rect 4692 -5966 4698 -5906
rect 4758 -5966 4764 -5906
rect 4562 -6078 4568 -6018
rect 4628 -6078 4634 -6018
rect 4698 -6154 4758 -5966
rect 4702 -7190 4762 -6856
rect 5208 -6940 5268 -6710
rect 5722 -6940 5782 -6856
rect 6228 -6940 6288 -6750
rect 5202 -7000 5208 -6940
rect 5268 -7000 6288 -6940
rect 5208 -7308 5268 -7000
rect 5722 -7194 5782 -7000
rect 6228 -7288 6288 -7000
rect 6360 -7050 6420 -5020
rect 6354 -7110 6360 -7050
rect 6420 -7110 6426 -7050
rect 4582 -8074 4642 -7888
rect 4694 -8034 4700 -7974
rect 4760 -8034 4766 -7974
rect 6360 -8028 6420 -7110
rect 6546 -7238 6552 -7178
rect 6612 -7238 6618 -7178
rect 4576 -8134 4582 -8074
rect 4642 -8134 4648 -8074
rect 4700 -8224 4760 -8034
rect 5208 -8088 6420 -8028
rect 5208 -8314 5268 -8088
rect 5710 -8226 5770 -8088
rect 6228 -8352 6288 -8088
rect 1402 -9084 1462 -9078
rect 3682 -9084 3742 -8916
rect 1462 -9144 3742 -9084
rect 1402 -9150 1462 -9144
rect 1542 -9260 1602 -9254
rect 4688 -9260 4748 -8909
rect 1602 -9320 4748 -9260
rect 1542 -9326 1602 -9320
rect 2442 -9434 2502 -9428
rect 5210 -9434 5270 -8778
rect 2502 -9494 5270 -9434
rect 2442 -9500 2502 -9494
rect 1282 -9584 1342 -9578
rect 6552 -9584 6612 -7238
rect 6686 -8330 6746 -4402
rect 6796 -5012 6802 -4952
rect 6862 -5012 6868 -4952
rect 6802 -7074 6862 -5012
rect 7044 -5916 7104 -1654
rect 7488 -1784 7552 -1654
rect 7482 -1848 7488 -1784
rect 7552 -1848 7558 -1784
rect 7312 -1934 7372 -1928
rect 7312 -4870 7372 -1994
rect 7990 -2040 8050 -1446
rect 8510 -1536 8570 -1350
rect 10546 -1362 10606 -1360
rect 8504 -1596 8510 -1536
rect 8570 -1596 8576 -1536
rect 9032 -2040 9092 -1440
rect 9526 -1646 9590 -1362
rect 9520 -1710 9526 -1646
rect 9590 -1710 9596 -1646
rect 10032 -2040 10092 -1446
rect 10546 -1536 10610 -1362
rect 11068 -1536 11128 -1436
rect 11566 -1536 11626 -1330
rect 12580 -1354 12640 -1352
rect 10540 -1596 10546 -1536
rect 10606 -1596 10612 -1536
rect 11062 -1596 11068 -1536
rect 11128 -1596 11134 -1536
rect 11560 -1596 11566 -1536
rect 11626 -1596 11632 -1536
rect 12040 -1540 12100 -1444
rect 12580 -1532 12644 -1354
rect 7422 -2100 7428 -2040
rect 7488 -2100 7494 -2040
rect 7984 -2100 7990 -2040
rect 8050 -2100 8056 -2040
rect 9026 -2100 9032 -2040
rect 9092 -2100 9098 -2040
rect 10026 -2100 10032 -2040
rect 10092 -2100 10098 -2040
rect 7428 -4682 7488 -2100
rect 12040 -2138 12100 -1600
rect 12548 -1536 12644 -1532
rect 12548 -1538 12580 -1536
rect 12640 -1596 12646 -1536
rect 13034 -1596 13040 -1536
rect 13100 -1596 13106 -1536
rect 12548 -2138 12608 -1598
rect 13040 -2138 13100 -1596
rect 13194 -2040 13254 -1444
rect 13598 -1788 13662 -1354
rect 13598 -1858 13662 -1852
rect 14084 -1534 14144 -1528
rect 13188 -2100 13194 -2040
rect 13254 -2100 13260 -2040
rect 14084 -2138 14144 -1594
rect 14204 -2040 14264 -1444
rect 14616 -1536 14676 -1326
rect 16654 -1346 16714 -1344
rect 14610 -1596 14616 -1536
rect 14676 -1596 14682 -1536
rect 15146 -2040 15206 -1444
rect 15634 -1930 15698 -1350
rect 16128 -1534 16188 -1528
rect 16654 -1534 16718 -1346
rect 15628 -1994 15634 -1930
rect 15698 -1994 15704 -1930
rect 14198 -2100 14204 -2040
rect 14264 -2100 14270 -2040
rect 15140 -2100 15146 -2040
rect 15206 -2100 15212 -2040
rect 16128 -2138 16188 -1594
rect 16622 -1538 16718 -1534
rect 16622 -1540 16654 -1538
rect 16714 -1598 16720 -1538
rect 17150 -1544 17210 -1430
rect 17672 -1534 17732 -940
rect 18690 -1358 18750 -1356
rect 16622 -2138 16682 -1600
rect 17150 -2138 17210 -1604
rect 17638 -1540 17732 -1534
rect 17698 -1542 17732 -1540
rect 17638 -1602 17672 -1600
rect 17638 -1608 17732 -1602
rect 18150 -1544 18210 -1436
rect 18690 -1540 18754 -1358
rect 18684 -1600 18690 -1540
rect 18750 -1600 18756 -1540
rect 17638 -2138 17698 -1608
rect 18150 -2138 18210 -1604
rect 19706 -1646 19770 -1352
rect 20724 -1358 20784 -1356
rect 20724 -1540 20788 -1358
rect 20718 -1600 20724 -1540
rect 20784 -1600 20790 -1540
rect 19700 -1710 19706 -1646
rect 19770 -1710 19776 -1646
rect 21740 -1934 21800 -1298
rect 22996 -1778 23056 680
rect 22992 -1784 23056 -1778
rect 22992 -1854 23056 -1848
rect 21734 -1994 21740 -1934
rect 21800 -1994 21806 -1934
rect 9704 -2198 19944 -2138
rect 7536 -2302 7542 -2242
rect 7602 -2302 7608 -2242
rect 7542 -4216 7602 -2302
rect 7668 -3176 7728 -2994
rect 8180 -3176 8240 -3086
rect 8686 -3176 8746 -3000
rect 7668 -3178 8746 -3176
rect 7668 -3236 8686 -3178
rect 8680 -3238 8686 -3236
rect 8746 -3238 8752 -3178
rect 9190 -3286 9250 -3084
rect 9184 -3346 9190 -3286
rect 9250 -3346 9256 -3286
rect 9190 -3424 9250 -3346
rect 7668 -4216 7728 -4000
rect 8170 -4216 8230 -4110
rect 8682 -4210 8742 -4026
rect 8676 -4216 8682 -4210
rect 7542 -4270 8682 -4216
rect 8742 -4270 8748 -4210
rect 7542 -4276 8748 -4270
rect 9188 -4344 9248 -4122
rect 9188 -4410 9248 -4404
rect 9704 -4552 9764 -2198
rect 10714 -2302 10720 -2242
rect 10780 -2302 10786 -2242
rect 10720 -2512 10780 -2302
rect 10210 -3280 10270 -3071
rect 10714 -3238 10720 -3178
rect 10780 -3238 10786 -3178
rect 10210 -3286 10272 -3280
rect 10210 -3346 10212 -3286
rect 10210 -3352 10272 -3346
rect 10210 -3414 10270 -3352
rect 10720 -3526 10780 -3238
rect 11232 -3280 11292 -3091
rect 11230 -3286 11292 -3280
rect 11290 -3346 11292 -3286
rect 11230 -3352 11292 -3346
rect 11232 -3434 11292 -3352
rect 10202 -4348 10262 -4106
rect 11234 -4340 11294 -4118
rect 11234 -4406 11294 -4400
rect 10202 -4414 10262 -4408
rect 11742 -4552 11802 -2198
rect 12252 -3280 12312 -3081
rect 12762 -3178 12822 -2960
rect 12756 -3238 12762 -3178
rect 12822 -3238 12828 -3178
rect 12252 -3286 12314 -3280
rect 12252 -3346 12254 -3286
rect 12252 -3352 12314 -3346
rect 13268 -3286 13328 -3075
rect 12252 -3424 12312 -3352
rect 13268 -3418 13328 -3346
rect 12232 -4340 12292 -4112
rect 12762 -4210 12822 -3990
rect 12756 -4270 12762 -4210
rect 12822 -4270 12828 -4210
rect 12232 -4406 12292 -4400
rect 13276 -4340 13336 -4096
rect 13276 -4406 13336 -4400
rect 13780 -4552 13840 -2198
rect 14782 -2302 14788 -2242
rect 14848 -2302 14854 -2242
rect 14788 -2522 14848 -2302
rect 14284 -3280 14344 -3081
rect 14782 -3238 14788 -3178
rect 14848 -3238 14854 -3178
rect 14284 -3286 14346 -3280
rect 14284 -3346 14286 -3286
rect 14284 -3352 14346 -3346
rect 14284 -3424 14344 -3352
rect 14788 -3542 14848 -3238
rect 15294 -3280 15354 -3081
rect 15294 -3286 15356 -3280
rect 15294 -3346 15296 -3286
rect 15294 -3352 15356 -3346
rect 15294 -3424 15354 -3352
rect 14280 -4344 14340 -4106
rect 14280 -4410 14340 -4404
rect 14798 -4460 14858 -3964
rect 15296 -4344 15356 -4102
rect 15296 -4410 15356 -4404
rect 14588 -4520 14858 -4460
rect 9704 -4612 14080 -4552
rect 14140 -4612 14146 -4552
rect 7428 -4742 11596 -4682
rect 7306 -4930 7312 -4870
rect 7372 -4930 7378 -4870
rect 8472 -4930 8478 -4870
rect 8538 -4930 8544 -4870
rect 7038 -5976 7044 -5916
rect 7104 -5976 7110 -5916
rect 6796 -7134 6802 -7074
rect 6862 -7134 6868 -7074
rect 6792 -7348 6798 -7288
rect 6858 -7348 6864 -7288
rect 6680 -8390 6686 -8330
rect 6746 -8390 6752 -8330
rect 1342 -9644 6612 -9584
rect 1282 -9650 1342 -9644
rect -13992 -10378 -2722 -10122
rect 372 -10242 484 -9728
rect 2336 -9846 2396 -9840
rect 6798 -9846 6858 -7348
rect 7044 -9588 7104 -5976
rect 7174 -6074 7180 -6014
rect 7240 -6074 7246 -6014
rect 7038 -9648 7044 -9588
rect 7104 -9648 7110 -9588
rect 7180 -9718 7240 -6074
rect 7312 -8538 7372 -4930
rect 8478 -5110 8538 -4930
rect 9494 -5130 9554 -4742
rect 10508 -4930 10514 -4870
rect 10574 -4930 10580 -4870
rect 10514 -5108 10574 -4930
rect 11016 -4934 11022 -4870
rect 11086 -4934 11092 -4870
rect 11022 -5028 11086 -4934
rect 11536 -5138 11596 -4742
rect 12040 -5028 12100 -4612
rect 7460 -5818 7520 -5624
rect 7974 -5818 8034 -5722
rect 8476 -5818 8536 -5636
rect 7460 -5878 8536 -5818
rect 8966 -6120 9026 -5714
rect 9496 -5818 9556 -5636
rect 9490 -5878 9496 -5818
rect 9556 -5878 9562 -5818
rect 10004 -5872 10064 -5713
rect 11010 -5872 11070 -5713
rect 11532 -5818 11592 -5632
rect 12042 -5814 12102 -5718
rect 12548 -5814 12608 -4612
rect 13040 -5024 13100 -4612
rect 14078 -5022 14138 -4612
rect 13062 -5814 13122 -5722
rect 13568 -5814 13628 -5636
rect 14072 -5814 14132 -5720
rect 9496 -6014 9556 -5878
rect 10004 -5932 11070 -5872
rect 11526 -5878 11532 -5818
rect 11592 -5878 11598 -5818
rect 11868 -5876 11874 -5816
rect 11934 -5876 11940 -5816
rect 12042 -5874 14132 -5814
rect 14588 -5816 14648 -4520
rect 15816 -4552 15876 -2198
rect 17846 -2858 17906 -2198
rect 18858 -2302 18864 -2242
rect 18924 -2302 18930 -2242
rect 18864 -2512 18924 -2302
rect 16316 -3280 16376 -3075
rect 16830 -3178 16890 -2960
rect 16824 -3238 16830 -3178
rect 16890 -3238 16896 -3178
rect 17330 -3280 17390 -3075
rect 16316 -3286 16378 -3280
rect 16316 -3346 16318 -3286
rect 16316 -3352 16378 -3346
rect 17330 -3286 17392 -3280
rect 17330 -3346 17332 -3286
rect 17330 -3352 17392 -3346
rect 16316 -3418 16376 -3352
rect 17330 -3418 17390 -3352
rect 16300 -4344 16360 -4112
rect 16830 -4210 16890 -3974
rect 16824 -4270 16830 -4210
rect 16890 -4270 16896 -4210
rect 16300 -4410 16360 -4404
rect 17332 -4340 17392 -4118
rect 17332 -4406 17392 -4400
rect 15090 -4812 15096 -4748
rect 15160 -4812 15166 -4748
rect 15096 -4870 15160 -4812
rect 15816 -4842 15876 -4612
rect 17846 -4452 17906 -2952
rect 18362 -3280 18422 -3075
rect 18860 -3238 18866 -3178
rect 18926 -3238 18932 -3178
rect 18362 -3286 18424 -3280
rect 18362 -3346 18364 -3286
rect 18362 -3352 18424 -3346
rect 18362 -3418 18422 -3352
rect 18866 -3548 18926 -3238
rect 19372 -3280 19432 -3075
rect 19372 -3286 19434 -3280
rect 19372 -3346 19374 -3286
rect 19372 -3352 19434 -3346
rect 19372 -3418 19432 -3352
rect 18348 -4344 18408 -4106
rect 18348 -4410 18408 -4404
rect 19376 -4344 19436 -4112
rect 19376 -4410 19436 -4404
rect 19884 -4452 19944 -2198
rect 22054 -2302 22060 -2242
rect 22120 -2302 22126 -2242
rect 20394 -3280 20454 -3081
rect 20902 -3176 20962 -2948
rect 21424 -3176 21484 -3088
rect 21918 -3176 21978 -2998
rect 20902 -3178 21978 -3176
rect 20896 -3238 20902 -3178
rect 20962 -3236 21978 -3178
rect 20962 -3238 20968 -3236
rect 20394 -3286 20456 -3280
rect 20394 -3346 20396 -3286
rect 20394 -3352 20456 -3346
rect 20394 -3424 20454 -3352
rect 20396 -4344 20456 -4106
rect 20898 -4206 20958 -3980
rect 21386 -4206 21446 -4112
rect 21918 -4206 21978 -3984
rect 22060 -4206 22120 -2302
rect 20896 -4210 22120 -4206
rect 20892 -4270 20898 -4210
rect 20958 -4266 22120 -4210
rect 20958 -4270 20964 -4266
rect 22848 -4402 22854 -4342
rect 22914 -4402 22920 -4342
rect 20396 -4410 20456 -4404
rect 17846 -4512 19944 -4452
rect 17846 -4842 17906 -4512
rect 21708 -4628 21714 -4568
rect 21774 -4628 21780 -4568
rect 19154 -4812 19160 -4748
rect 19224 -4812 19230 -4748
rect 20178 -4812 20184 -4748
rect 20248 -4812 20254 -4748
rect 21190 -4812 21196 -4748
rect 21260 -4812 21266 -4748
rect 15092 -4934 15098 -4870
rect 15162 -4934 15168 -4870
rect 15816 -4902 18210 -4842
rect 19160 -4866 19224 -4812
rect 15096 -5022 15160 -4934
rect 16128 -5028 16188 -4902
rect 9490 -6074 9496 -6014
rect 9556 -6074 9562 -6014
rect 10004 -6120 10064 -5932
rect 10510 -6072 10516 -6012
rect 10576 -6072 10582 -6012
rect 8476 -6184 8482 -6124
rect 8542 -6184 8548 -6124
rect 8966 -6180 10064 -6120
rect 10516 -6124 10576 -6072
rect 8482 -6366 8542 -6184
rect 8966 -6282 9026 -6180
rect 10004 -6287 10064 -6180
rect 10510 -6184 10516 -6124
rect 10576 -6184 10582 -6124
rect 10516 -6362 10576 -6184
rect 11010 -6287 11070 -5932
rect 11874 -6130 11934 -5876
rect 11532 -6190 11934 -6130
rect 11532 -6398 11592 -6190
rect 12548 -6384 12608 -5874
rect 14582 -5876 14588 -5816
rect 14648 -5876 14654 -5816
rect 15606 -6012 15666 -5582
rect 16116 -5814 16176 -5722
rect 16622 -5814 16682 -4902
rect 17150 -5032 17210 -4902
rect 17142 -5814 17202 -5721
rect 17638 -5814 17698 -4902
rect 18150 -5038 18210 -4902
rect 18654 -4930 18660 -4870
rect 18720 -4930 18726 -4870
rect 18660 -5112 18720 -4930
rect 19160 -5028 19224 -4930
rect 20184 -5022 20248 -4812
rect 20688 -4930 20694 -4870
rect 20754 -4930 20760 -4870
rect 20694 -5108 20754 -4930
rect 21196 -5018 21260 -4812
rect 21714 -4866 21774 -4628
rect 21714 -4926 22790 -4866
rect 21714 -5120 21774 -4926
rect 22228 -5022 22288 -4926
rect 22730 -5108 22790 -4926
rect 18154 -5814 18214 -5724
rect 16116 -5874 18214 -5814
rect 15600 -6072 15606 -6012
rect 15666 -6072 15672 -6012
rect 13566 -6186 13572 -6126
rect 13632 -6186 13638 -6126
rect 15600 -6186 15606 -6126
rect 15666 -6186 15672 -6126
rect 13572 -6368 13632 -6186
rect 15606 -6370 15666 -6186
rect 17638 -6360 17698 -5874
rect 18656 -6186 18662 -6126
rect 18722 -6186 18728 -6126
rect 18662 -6368 18722 -6186
rect 19162 -6287 19222 -5713
rect 19676 -5818 19736 -5636
rect 19670 -5878 19676 -5818
rect 19736 -5878 19742 -5818
rect 20186 -6287 20246 -5713
rect 20690 -6186 20696 -6126
rect 20756 -6186 20762 -6126
rect 20696 -6364 20756 -6186
rect 21192 -6281 21252 -5707
rect 21712 -5818 21772 -5632
rect 21706 -5878 21712 -5818
rect 21772 -5878 21778 -5818
rect 21714 -6180 22790 -6120
rect 21714 -6374 21774 -6180
rect 22228 -6276 22288 -6180
rect 22730 -6362 22790 -6180
rect 7464 -7074 7524 -6880
rect 7978 -7074 8038 -6978
rect 8480 -7074 8540 -6892
rect 7464 -7134 8540 -7074
rect 7464 -7288 7524 -7134
rect 7458 -7348 7464 -7288
rect 7524 -7348 7530 -7288
rect 7462 -7458 8538 -7398
rect 7462 -7630 7522 -7458
rect 7976 -7532 8036 -7458
rect 8478 -7618 8538 -7458
rect 8960 -7542 9020 -6968
rect 9498 -7178 9558 -6890
rect 9498 -7244 9558 -7238
rect 9492 -7442 9498 -7382
rect 9558 -7442 9564 -7382
rect 9498 -7620 9558 -7442
rect 9998 -7543 10058 -6968
rect 11004 -7543 11064 -6968
rect 11534 -7178 11594 -6886
rect 12054 -7070 12114 -6977
rect 12550 -7070 12610 -6886
rect 13066 -7070 13126 -6980
rect 12054 -7130 13126 -7070
rect 11528 -7238 11534 -7178
rect 11594 -7238 11600 -7178
rect 11526 -7340 11532 -7280
rect 11592 -7340 11598 -7280
rect 11532 -7382 11592 -7340
rect 11526 -7442 11532 -7382
rect 11592 -7442 11598 -7382
rect 11532 -7624 11592 -7442
rect 12550 -7634 12610 -7130
rect 13562 -7134 13568 -7074
rect 13628 -7134 13634 -7074
rect 13568 -7620 13628 -7134
rect 14070 -7236 14130 -6974
rect 14588 -7074 14648 -6892
rect 14582 -7134 14588 -7074
rect 14648 -7134 14654 -7074
rect 15100 -7236 15160 -6962
rect 14070 -7296 15160 -7236
rect 14070 -7548 14130 -7296
rect 14582 -7440 14588 -7380
rect 14648 -7440 14654 -7380
rect 14588 -7618 14648 -7440
rect 15100 -7536 15160 -7296
rect 15606 -7380 15666 -6888
rect 15600 -7440 15606 -7380
rect 15666 -7440 15672 -7380
rect 16112 -7536 16172 -6962
rect 16624 -7074 16684 -6888
rect 17142 -7072 17202 -6979
rect 17638 -7072 17698 -6888
rect 18154 -7072 18214 -6982
rect 16618 -7134 16624 -7074
rect 16684 -7134 16690 -7074
rect 17142 -7132 18214 -7072
rect 16616 -7440 16622 -7380
rect 16682 -7440 16688 -7380
rect 16622 -7622 16682 -7440
rect 17638 -7626 17698 -7132
rect 18652 -7238 18658 -7178
rect 18718 -7238 18724 -7178
rect 18658 -7628 18718 -7238
rect 19156 -7543 19216 -6968
rect 19520 -7120 19526 -7060
rect 19586 -7120 19592 -7060
rect 19526 -7380 19586 -7120
rect 19674 -7170 19734 -6880
rect 19668 -7230 19674 -7170
rect 19734 -7230 19740 -7170
rect 19520 -7440 19526 -7380
rect 19586 -7440 19592 -7380
rect 19672 -7438 19678 -7378
rect 19738 -7438 19744 -7378
rect 19678 -7616 19738 -7438
rect 20180 -7543 20240 -6968
rect 20694 -7280 20754 -6888
rect 20688 -7340 20694 -7280
rect 20754 -7340 20760 -7280
rect 21186 -7537 21246 -6962
rect 21714 -7170 21774 -6876
rect 22854 -7170 22914 -4402
rect 22996 -4570 23056 -1854
rect 23284 -4270 23290 -4210
rect 23350 -4270 23356 -4210
rect 22996 -4636 23056 -4630
rect 23132 -4930 23138 -4870
rect 23198 -4930 23204 -4870
rect 22972 -6072 22978 -6012
rect 23038 -6072 23044 -6012
rect 21708 -7230 21714 -7170
rect 21774 -7230 21780 -7170
rect 22848 -7230 22854 -7170
rect 22914 -7230 22920 -7170
rect 21706 -7438 21712 -7378
rect 21772 -7438 21778 -7378
rect 21712 -7620 21772 -7438
rect 8480 -8330 8540 -8144
rect 8474 -8390 8480 -8330
rect 8540 -8390 8546 -8330
rect 7306 -8598 7312 -8538
rect 7372 -8598 7378 -8538
rect 7462 -8696 8538 -8636
rect 7462 -8890 7522 -8696
rect 7976 -8792 8036 -8696
rect 8478 -8878 8538 -8696
rect 8972 -8792 9032 -8218
rect 9488 -8700 9494 -8640
rect 9554 -8700 9560 -8640
rect 9494 -8878 9554 -8700
rect 10010 -8792 10070 -8218
rect 10516 -8330 10576 -8148
rect 10510 -8390 10516 -8330
rect 10576 -8390 10582 -8330
rect 10516 -8438 10576 -8390
rect 10510 -8498 10516 -8438
rect 10576 -8498 10582 -8438
rect 11016 -8488 11076 -8218
rect 11534 -8322 11594 -8153
rect 12052 -8322 12112 -8229
rect 12548 -8322 12608 -8138
rect 13064 -8322 13124 -8232
rect 11528 -8382 11534 -8322
rect 11594 -8382 11600 -8322
rect 12052 -8382 13124 -8322
rect 13330 -8382 13336 -8322
rect 13396 -8382 13402 -8322
rect 13570 -8328 13630 -8142
rect 11016 -8548 11792 -8488
rect 11016 -8792 11076 -8548
rect 11522 -8700 11528 -8640
rect 11588 -8700 11594 -8640
rect 11732 -8652 11792 -8548
rect 11528 -8882 11588 -8700
rect 11726 -8712 11732 -8652
rect 11792 -8712 11798 -8652
rect 12548 -8910 12608 -8382
rect 13336 -8592 13396 -8382
rect 13564 -8388 13570 -8328
rect 13630 -8388 13636 -8328
rect 14066 -8450 14126 -8228
rect 15094 -8450 15154 -8234
rect 15606 -8328 15666 -8146
rect 15600 -8388 15606 -8328
rect 15666 -8388 15672 -8328
rect 14066 -8510 15154 -8450
rect 15598 -8498 15604 -8438
rect 15664 -8498 15670 -8438
rect 13336 -8652 14644 -8592
rect 14584 -8904 14644 -8652
rect 15094 -8652 15154 -8510
rect 15094 -8790 15154 -8712
rect 15604 -8916 15664 -8498
rect 16110 -8652 16170 -8226
rect 17140 -8324 17200 -8231
rect 17636 -8324 17696 -8140
rect 18152 -8324 18212 -8234
rect 17140 -8384 18212 -8324
rect 18660 -8326 18720 -8140
rect 16110 -8718 16170 -8712
rect 17636 -8890 17696 -8384
rect 18654 -8386 18660 -8326
rect 18720 -8386 18726 -8326
rect 19168 -8646 19228 -8218
rect 19168 -8652 19230 -8646
rect 19168 -8712 19170 -8652
rect 19676 -8700 19682 -8640
rect 19742 -8700 19748 -8640
rect 19168 -8718 19230 -8712
rect 19168 -8792 19228 -8718
rect 19682 -8878 19742 -8700
rect 20192 -8792 20252 -8218
rect 20696 -8326 20756 -8144
rect 20690 -8386 20696 -8326
rect 20756 -8386 20762 -8326
rect 21198 -8786 21258 -8212
rect 21712 -8330 21772 -8136
rect 22226 -8330 22286 -8234
rect 22728 -8330 22788 -8148
rect 21712 -8390 22788 -8330
rect 22854 -8438 22914 -7230
rect 22978 -7378 23038 -6072
rect 22972 -7438 22978 -7378
rect 23038 -7438 23044 -7378
rect 22848 -8498 22854 -8438
rect 22914 -8498 22920 -8438
rect 21710 -8700 21716 -8640
rect 21776 -8700 21782 -8640
rect 21716 -8882 21776 -8700
rect 8476 -9588 8536 -9402
rect 8470 -9648 8476 -9588
rect 8536 -9648 8542 -9588
rect 8984 -9702 9044 -9490
rect 10008 -9702 10068 -9482
rect 10512 -9588 10572 -9406
rect 10506 -9648 10512 -9588
rect 10572 -9648 10578 -9588
rect 11014 -9702 11074 -9482
rect 7174 -9778 7180 -9718
rect 7240 -9778 7246 -9718
rect 8984 -9762 11074 -9702
rect 2332 -9906 2336 -9846
rect 2396 -9906 6858 -9846
rect 2336 -9912 2396 -9906
rect 2216 -9964 2276 -9958
rect 7180 -9964 7240 -9778
rect 2276 -10024 7240 -9964
rect 2216 -10030 2276 -10024
rect 1770 -10082 1830 -10076
rect 8984 -10082 9044 -9762
rect 11014 -9972 11074 -9762
rect 11534 -9858 11594 -9392
rect 12052 -9582 12112 -9487
rect 12548 -9582 12608 -9396
rect 13064 -9582 13124 -9490
rect 13570 -9582 13630 -9384
rect 14080 -9582 14140 -9490
rect 16106 -9582 16166 -9490
rect 16622 -9582 16682 -9400
rect 17140 -9582 17200 -9489
rect 17636 -9582 17696 -9398
rect 18152 -9582 18212 -9492
rect 12052 -9642 18212 -9582
rect 18664 -9588 18724 -9402
rect 18658 -9648 18664 -9588
rect 18724 -9648 18730 -9588
rect 19172 -9700 19232 -9474
rect 20192 -9700 20252 -9482
rect 20700 -9588 20760 -9406
rect 20694 -9648 20700 -9588
rect 20760 -9648 20766 -9588
rect 21194 -9700 21254 -9482
rect 21714 -9584 21774 -9390
rect 22228 -9584 22288 -9488
rect 22730 -9584 22790 -9402
rect 21714 -9644 22790 -9584
rect 19172 -9760 21254 -9700
rect 11528 -9918 11534 -9858
rect 11594 -9918 11600 -9858
rect 19172 -9972 19232 -9760
rect 23138 -9858 23198 -4930
rect 23290 -6126 23350 -4270
rect 23284 -6186 23290 -6126
rect 23350 -6186 23356 -6126
rect 24716 -9728 24722 3702
rect 24822 -9728 24828 3702
rect 23132 -9918 23138 -9858
rect 23198 -9918 23204 -9858
rect 11014 -10032 19232 -9972
rect 1830 -10142 9044 -10082
rect 1770 -10148 1830 -10142
rect 24716 -10242 24828 -9728
rect 372 -10248 24828 -10242
rect 372 -10348 478 -10248
rect 24722 -10348 24828 -10248
rect 372 -10354 24828 -10348
rect -13992 -10670 -13630 -10378
rect -2866 -10670 -2722 -10378
rect -13992 -10978 -2722 -10670
rect -13992 -11172 -1640 -10978
rect -13992 -11178 24928 -11172
rect -13992 -11278 -12222 -11178
rect 24822 -11278 24928 -11178
rect -13992 -11284 24928 -11278
rect -13992 -11300 -1642 -11284
rect -12328 -12070 -12216 -11300
rect 1888 -11358 1948 -11352
rect 2210 -11408 2216 -11348
rect 2276 -11408 2282 -11348
rect 2336 -11356 2396 -11350
rect 1276 -11554 1282 -11494
rect 1342 -11554 1348 -11494
rect 1396 -11552 1402 -11492
rect 1462 -11552 1468 -11492
rect 1536 -11534 1542 -11474
rect 1602 -11534 1608 -11474
rect 1764 -11518 1770 -11458
rect 1830 -11518 1836 -11458
rect 1144 -11682 1150 -11622
rect 1210 -11682 1216 -11622
rect -12328 -26330 -12322 -12070
rect -12222 -26330 -12216 -12070
rect -1568 -12280 -1562 -12220
rect -1502 -12280 -1496 -12220
rect -1562 -12324 -1502 -12280
rect -9196 -12384 -1502 -12324
rect -9196 -12524 -9136 -12384
rect -8686 -12434 -8626 -12384
rect -8902 -12440 -8414 -12434
rect -8902 -12474 -8890 -12440
rect -8426 -12474 -8414 -12440
rect -8902 -12480 -8414 -12474
rect -9196 -12554 -9184 -12524
rect -9190 -13082 -9184 -12554
rect -9200 -13100 -9184 -13082
rect -9150 -12554 -9136 -12524
rect -8180 -12524 -8120 -12384
rect -7678 -12434 -7618 -12384
rect -6650 -12434 -6590 -12384
rect -7884 -12440 -7396 -12434
rect -7884 -12474 -7872 -12440
rect -7408 -12474 -7396 -12440
rect -7884 -12480 -7396 -12474
rect -6866 -12440 -6378 -12434
rect -6866 -12474 -6854 -12440
rect -6390 -12474 -6378 -12440
rect -6866 -12480 -6378 -12474
rect -8180 -12548 -8166 -12524
rect -9150 -13082 -9144 -12554
rect -8172 -13078 -8166 -12548
rect -9150 -13100 -9140 -13082
rect -9200 -13342 -9140 -13100
rect -8180 -13100 -8166 -13078
rect -8132 -12548 -8120 -12524
rect -7154 -12524 -7108 -12512
rect -8132 -13078 -8126 -12548
rect -7154 -13076 -7148 -12524
rect -8132 -13100 -8120 -13078
rect -8902 -13150 -8414 -13144
rect -8902 -13184 -8890 -13150
rect -8426 -13184 -8414 -13150
rect -8902 -13190 -8414 -13184
rect -8686 -13252 -8626 -13190
rect -8902 -13258 -8414 -13252
rect -8902 -13292 -8890 -13258
rect -8426 -13292 -8414 -13258
rect -8902 -13298 -8414 -13292
rect -9200 -13372 -9184 -13342
rect -9190 -13896 -9184 -13372
rect -9198 -13918 -9184 -13896
rect -9150 -13372 -9140 -13342
rect -8180 -13342 -8120 -13100
rect -7160 -13100 -7148 -13076
rect -7114 -13076 -7108 -12524
rect -6142 -12524 -6082 -12384
rect -5636 -12434 -5576 -12384
rect -4622 -12434 -4562 -12384
rect -5848 -12440 -5360 -12434
rect -5848 -12474 -5836 -12440
rect -5372 -12474 -5360 -12440
rect -5848 -12480 -5360 -12474
rect -4830 -12440 -4342 -12434
rect -4830 -12474 -4818 -12440
rect -4354 -12474 -4342 -12440
rect -4830 -12480 -4342 -12474
rect -6142 -12562 -6130 -12524
rect -7114 -13100 -7100 -13076
rect -6136 -13080 -6130 -12562
rect -7884 -13150 -7396 -13144
rect -7884 -13184 -7872 -13150
rect -7408 -13184 -7396 -13150
rect -7884 -13190 -7396 -13184
rect -7682 -13252 -7622 -13190
rect -7884 -13258 -7396 -13252
rect -7884 -13292 -7872 -13258
rect -7408 -13292 -7396 -13258
rect -7884 -13298 -7396 -13292
rect -8180 -13368 -8166 -13342
rect -9150 -13896 -9144 -13372
rect -8172 -13892 -8166 -13368
rect -9150 -13918 -9138 -13896
rect -9198 -14160 -9138 -13918
rect -8178 -13918 -8166 -13892
rect -8132 -13368 -8120 -13342
rect -7160 -13342 -7100 -13100
rect -6142 -13100 -6130 -13080
rect -6096 -12562 -6082 -12524
rect -5118 -12524 -5072 -12512
rect -4106 -12524 -4046 -12384
rect -3590 -12434 -3530 -12384
rect -2584 -12434 -2524 -12384
rect -3812 -12440 -3324 -12434
rect -3812 -12474 -3800 -12440
rect -3336 -12474 -3324 -12440
rect -3812 -12480 -3324 -12474
rect -2794 -12440 -2306 -12434
rect -2794 -12474 -2782 -12440
rect -2318 -12474 -2306 -12440
rect -2794 -12480 -2306 -12474
rect -6096 -13080 -6090 -12562
rect -5118 -13072 -5112 -12524
rect -6096 -13100 -6082 -13080
rect -6866 -13150 -6378 -13144
rect -6866 -13184 -6854 -13150
rect -6390 -13184 -6378 -13150
rect -6866 -13190 -6378 -13184
rect -6652 -13252 -6592 -13190
rect -6866 -13258 -6378 -13252
rect -6866 -13292 -6854 -13258
rect -6390 -13292 -6378 -13258
rect -6866 -13298 -6378 -13292
rect -7160 -13366 -7148 -13342
rect -8132 -13892 -8126 -13368
rect -7154 -13890 -7148 -13366
rect -8132 -13918 -8118 -13892
rect -8902 -13968 -8414 -13962
rect -8902 -14002 -8890 -13968
rect -8426 -14002 -8414 -13968
rect -8902 -14008 -8414 -14002
rect -8686 -14070 -8626 -14008
rect -8902 -14076 -8414 -14070
rect -8902 -14110 -8890 -14076
rect -8426 -14110 -8414 -14076
rect -8902 -14116 -8414 -14110
rect -9198 -14186 -9184 -14160
rect -9190 -14724 -9184 -14186
rect -9198 -14736 -9184 -14724
rect -9150 -14186 -9138 -14160
rect -8178 -14160 -8118 -13918
rect -7158 -13918 -7148 -13890
rect -7114 -13366 -7100 -13342
rect -6142 -13342 -6082 -13100
rect -5122 -13100 -5112 -13072
rect -5078 -13072 -5072 -12524
rect -4108 -12558 -4094 -12524
rect -4106 -12570 -4094 -12558
rect -5078 -13100 -5062 -13072
rect -4100 -13080 -4094 -12570
rect -5848 -13150 -5360 -13144
rect -5848 -13184 -5836 -13150
rect -5372 -13184 -5360 -13150
rect -5848 -13190 -5360 -13184
rect -5650 -13252 -5590 -13190
rect -5848 -13258 -5360 -13252
rect -5848 -13292 -5836 -13258
rect -5372 -13292 -5360 -13258
rect -5848 -13298 -5360 -13292
rect -7114 -13890 -7108 -13366
rect -6142 -13370 -6130 -13342
rect -7114 -13918 -7098 -13890
rect -6136 -13894 -6130 -13370
rect -7884 -13968 -7396 -13962
rect -7884 -14002 -7872 -13968
rect -7408 -14002 -7396 -13968
rect -7884 -14008 -7396 -14002
rect -7670 -14070 -7610 -14008
rect -7884 -14076 -7396 -14070
rect -7884 -14110 -7872 -14076
rect -7408 -14110 -7396 -14076
rect -7884 -14116 -7396 -14110
rect -8178 -14182 -8166 -14160
rect -9150 -14724 -9144 -14186
rect -8172 -14720 -8166 -14182
rect -9150 -14736 -9138 -14724
rect -9198 -14978 -9138 -14736
rect -8178 -14736 -8166 -14720
rect -8132 -14182 -8118 -14160
rect -7158 -14160 -7098 -13918
rect -6140 -13918 -6130 -13894
rect -6096 -13370 -6082 -13342
rect -5122 -13342 -5062 -13100
rect -4110 -13100 -4094 -13080
rect -4060 -12570 -4046 -12524
rect -3082 -12524 -3036 -12512
rect -4060 -13080 -4054 -12570
rect -3082 -13080 -3076 -12524
rect -4060 -13100 -4050 -13080
rect -4830 -13150 -4342 -13144
rect -4830 -13184 -4818 -13150
rect -4354 -13184 -4342 -13150
rect -4830 -13190 -4342 -13184
rect -4620 -13252 -4560 -13190
rect -4830 -13258 -4342 -13252
rect -4830 -13292 -4818 -13258
rect -4354 -13292 -4342 -13258
rect -4830 -13298 -4342 -13292
rect -5122 -13362 -5112 -13342
rect -6096 -13894 -6090 -13370
rect -5118 -13886 -5112 -13362
rect -6096 -13918 -6080 -13894
rect -6866 -13968 -6378 -13962
rect -6866 -14002 -6854 -13968
rect -6390 -14002 -6378 -13968
rect -6866 -14008 -6378 -14002
rect -6652 -14070 -6592 -14008
rect -6866 -14076 -6378 -14070
rect -6866 -14110 -6854 -14076
rect -6390 -14110 -6378 -14076
rect -6866 -14116 -6378 -14110
rect -7158 -14180 -7148 -14160
rect -8132 -14720 -8126 -14182
rect -7154 -14718 -7148 -14180
rect -8132 -14736 -8118 -14720
rect -8902 -14786 -8414 -14780
rect -8902 -14820 -8890 -14786
rect -8426 -14820 -8414 -14786
rect -8902 -14826 -8414 -14820
rect -8692 -14888 -8632 -14826
rect -8902 -14894 -8414 -14888
rect -8902 -14928 -8890 -14894
rect -8426 -14928 -8414 -14894
rect -8902 -14934 -8414 -14928
rect -9198 -15014 -9184 -14978
rect -9190 -15536 -9184 -15014
rect -9198 -15554 -9184 -15536
rect -9150 -15014 -9138 -14978
rect -8178 -14978 -8118 -14736
rect -7158 -14736 -7148 -14718
rect -7114 -14180 -7098 -14160
rect -6140 -14160 -6080 -13918
rect -5120 -13918 -5112 -13886
rect -5078 -13362 -5062 -13342
rect -4110 -13342 -4050 -13100
rect -3088 -13100 -3076 -13080
rect -3042 -13080 -3036 -12524
rect -2072 -12524 -2012 -12384
rect -1562 -12434 -1502 -12384
rect -42 -12414 -36 -12354
rect 24 -12414 30 -12354
rect -1776 -12440 -1288 -12434
rect -1776 -12474 -1764 -12440
rect -1300 -12474 -1288 -12440
rect -1776 -12480 -1288 -12474
rect -758 -12440 -270 -12434
rect -758 -12474 -746 -12440
rect -282 -12474 -270 -12440
rect -758 -12480 -270 -12474
rect -2072 -12560 -2058 -12524
rect -2064 -13080 -2058 -12560
rect -3042 -13100 -3028 -13080
rect -3812 -13150 -3324 -13144
rect -3812 -13184 -3800 -13150
rect -3336 -13184 -3324 -13150
rect -3812 -13190 -3324 -13184
rect -3604 -13252 -3544 -13190
rect -3812 -13258 -3324 -13252
rect -3812 -13292 -3800 -13258
rect -3336 -13292 -3324 -13258
rect -3812 -13298 -3324 -13292
rect -5078 -13886 -5072 -13362
rect -4110 -13370 -4094 -13342
rect -5078 -13918 -5060 -13886
rect -4100 -13894 -4094 -13370
rect -5848 -13968 -5360 -13962
rect -5848 -14002 -5836 -13968
rect -5372 -14002 -5360 -13968
rect -5848 -14008 -5360 -14002
rect -5650 -14070 -5590 -14008
rect -5848 -14076 -5360 -14070
rect -5848 -14110 -5836 -14076
rect -5372 -14110 -5360 -14076
rect -5848 -14116 -5360 -14110
rect -7114 -14718 -7108 -14180
rect -6140 -14184 -6130 -14160
rect -7114 -14736 -7098 -14718
rect -6136 -14722 -6130 -14184
rect -7884 -14786 -7396 -14780
rect -7884 -14820 -7872 -14786
rect -7408 -14820 -7396 -14786
rect -7884 -14826 -7396 -14820
rect -7670 -14888 -7610 -14826
rect -7884 -14894 -7396 -14888
rect -7884 -14928 -7872 -14894
rect -7408 -14928 -7396 -14894
rect -7884 -14934 -7396 -14928
rect -8178 -15010 -8166 -14978
rect -9150 -15536 -9144 -15014
rect -8172 -15532 -8166 -15010
rect -9150 -15554 -9138 -15536
rect -9198 -15796 -9138 -15554
rect -8178 -15554 -8166 -15532
rect -8132 -15010 -8118 -14978
rect -7158 -14978 -7098 -14736
rect -6140 -14736 -6130 -14722
rect -6096 -14184 -6080 -14160
rect -5120 -14160 -5060 -13918
rect -4108 -13918 -4094 -13894
rect -4060 -13370 -4050 -13342
rect -3088 -13342 -3028 -13100
rect -2068 -13100 -2058 -13080
rect -2024 -12560 -2012 -12524
rect -1046 -12524 -1000 -12512
rect -2024 -13080 -2018 -12560
rect -1046 -13076 -1040 -12524
rect -2024 -13100 -2008 -13080
rect -2794 -13150 -2306 -13144
rect -2794 -13184 -2782 -13150
rect -2318 -13184 -2306 -13150
rect -2794 -13190 -2306 -13184
rect -2582 -13252 -2522 -13190
rect -2794 -13258 -2306 -13252
rect -2794 -13292 -2782 -13258
rect -2318 -13292 -2306 -13258
rect -2794 -13298 -2306 -13292
rect -3088 -13370 -3076 -13342
rect -4060 -13894 -4054 -13370
rect -3082 -13894 -3076 -13370
rect -4060 -13918 -4048 -13894
rect -4830 -13968 -4342 -13962
rect -4830 -14002 -4818 -13968
rect -4354 -14002 -4342 -13968
rect -4830 -14008 -4342 -14002
rect -4620 -14070 -4560 -14008
rect -4830 -14076 -4342 -14070
rect -4830 -14110 -4818 -14076
rect -4354 -14110 -4342 -14076
rect -4830 -14116 -4342 -14110
rect -5120 -14176 -5112 -14160
rect -6096 -14722 -6090 -14184
rect -5118 -14714 -5112 -14176
rect -6096 -14736 -6080 -14722
rect -6866 -14786 -6378 -14780
rect -6866 -14820 -6854 -14786
rect -6390 -14820 -6378 -14786
rect -6866 -14826 -6378 -14820
rect -6658 -14888 -6598 -14826
rect -6866 -14894 -6378 -14888
rect -6866 -14928 -6854 -14894
rect -6390 -14928 -6378 -14894
rect -6866 -14934 -6378 -14928
rect -7158 -15008 -7148 -14978
rect -8132 -15532 -8126 -15010
rect -7154 -15530 -7148 -15008
rect -8132 -15554 -8118 -15532
rect -8902 -15604 -8414 -15598
rect -8902 -15638 -8890 -15604
rect -8426 -15638 -8414 -15604
rect -8902 -15644 -8414 -15638
rect -8694 -15706 -8634 -15644
rect -8902 -15712 -8414 -15706
rect -8902 -15746 -8890 -15712
rect -8426 -15746 -8414 -15712
rect -8902 -15752 -8414 -15746
rect -9198 -15826 -9184 -15796
rect -9190 -16356 -9184 -15826
rect -9198 -16372 -9184 -16356
rect -9150 -15826 -9138 -15796
rect -8178 -15796 -8118 -15554
rect -7158 -15554 -7148 -15530
rect -7114 -15008 -7098 -14978
rect -6140 -14978 -6080 -14736
rect -5120 -14736 -5112 -14714
rect -5078 -14176 -5060 -14160
rect -4108 -14160 -4048 -13918
rect -3086 -13918 -3076 -13894
rect -3042 -13370 -3028 -13342
rect -2068 -13342 -2008 -13100
rect -1052 -13100 -1040 -13076
rect -1006 -13076 -1000 -12524
rect -36 -12524 24 -12414
rect -36 -12560 -22 -12524
rect -1006 -13100 -992 -13076
rect -28 -13080 -22 -12560
rect -1776 -13150 -1288 -13144
rect -1776 -13184 -1764 -13150
rect -1300 -13184 -1288 -13150
rect -1776 -13190 -1288 -13184
rect -1570 -13252 -1510 -13190
rect -1776 -13258 -1288 -13252
rect -1776 -13292 -1764 -13258
rect -1300 -13292 -1288 -13258
rect -1776 -13298 -1288 -13292
rect -2068 -13370 -2058 -13342
rect -3042 -13894 -3036 -13370
rect -2064 -13894 -2058 -13370
rect -3042 -13918 -3026 -13894
rect -3812 -13968 -3324 -13962
rect -3812 -14002 -3800 -13968
rect -3336 -14002 -3324 -13968
rect -3812 -14008 -3324 -14002
rect -3604 -14070 -3544 -14008
rect -3812 -14076 -3324 -14070
rect -3812 -14110 -3800 -14076
rect -3336 -14110 -3324 -14076
rect -3812 -14116 -3324 -14110
rect -5078 -14714 -5072 -14176
rect -4108 -14184 -4094 -14160
rect -5078 -14736 -5060 -14714
rect -4100 -14722 -4094 -14184
rect -5848 -14786 -5360 -14780
rect -5848 -14820 -5836 -14786
rect -5372 -14820 -5360 -14786
rect -5848 -14826 -5360 -14820
rect -5656 -14888 -5596 -14826
rect -5848 -14894 -5360 -14888
rect -5848 -14928 -5836 -14894
rect -5372 -14928 -5360 -14894
rect -5848 -14934 -5360 -14928
rect -7114 -15530 -7108 -15008
rect -6140 -15012 -6130 -14978
rect -7114 -15554 -7098 -15530
rect -6136 -15534 -6130 -15012
rect -7884 -15604 -7396 -15598
rect -7884 -15638 -7872 -15604
rect -7408 -15638 -7396 -15604
rect -7884 -15644 -7396 -15638
rect -7676 -15706 -7616 -15644
rect -7884 -15712 -7396 -15706
rect -7884 -15746 -7872 -15712
rect -7408 -15746 -7396 -15712
rect -7884 -15752 -7396 -15746
rect -8178 -15822 -8166 -15796
rect -9150 -16356 -9144 -15826
rect -8172 -16352 -8166 -15822
rect -9150 -16372 -9138 -16356
rect -9198 -16614 -9138 -16372
rect -8178 -16372 -8166 -16352
rect -8132 -15822 -8118 -15796
rect -7158 -15796 -7098 -15554
rect -6140 -15554 -6130 -15534
rect -6096 -15012 -6080 -14978
rect -5120 -14978 -5060 -14736
rect -4108 -14736 -4094 -14722
rect -4060 -14184 -4048 -14160
rect -3086 -14160 -3026 -13918
rect -2066 -13918 -2058 -13894
rect -2024 -13370 -2008 -13342
rect -1052 -13342 -992 -13100
rect -30 -13100 -22 -13080
rect 12 -12560 24 -12524
rect 12 -13080 18 -12560
rect 12 -13100 30 -13080
rect -758 -13150 -270 -13144
rect -758 -13184 -746 -13150
rect -282 -13184 -270 -13150
rect -758 -13190 -270 -13184
rect -550 -13252 -490 -13190
rect -758 -13258 -270 -13252
rect -758 -13292 -746 -13258
rect -282 -13292 -270 -13258
rect -758 -13298 -270 -13292
rect -1052 -13366 -1040 -13342
rect -2024 -13894 -2018 -13370
rect -1046 -13890 -1040 -13366
rect -2024 -13918 -2006 -13894
rect -2794 -13968 -2306 -13962
rect -2794 -14002 -2782 -13968
rect -2318 -14002 -2306 -13968
rect -2794 -14008 -2306 -14002
rect -2582 -14070 -2522 -14008
rect -2794 -14076 -2306 -14070
rect -2794 -14110 -2782 -14076
rect -2318 -14110 -2306 -14076
rect -2794 -14116 -2306 -14110
rect -3086 -14184 -3076 -14160
rect -4060 -14722 -4054 -14184
rect -3082 -14722 -3076 -14184
rect -4060 -14736 -4048 -14722
rect -4830 -14786 -4342 -14780
rect -4830 -14820 -4818 -14786
rect -4354 -14820 -4342 -14786
rect -4830 -14826 -4342 -14820
rect -4626 -14888 -4566 -14826
rect -4830 -14894 -4342 -14888
rect -4830 -14928 -4818 -14894
rect -4354 -14928 -4342 -14894
rect -4830 -14934 -4342 -14928
rect -5120 -15004 -5112 -14978
rect -6096 -15534 -6090 -15012
rect -5118 -15526 -5112 -15004
rect -6096 -15554 -6080 -15534
rect -6866 -15604 -6378 -15598
rect -6866 -15638 -6854 -15604
rect -6390 -15638 -6378 -15604
rect -6866 -15644 -6378 -15638
rect -6660 -15706 -6600 -15644
rect -6866 -15712 -6378 -15706
rect -6866 -15746 -6854 -15712
rect -6390 -15746 -6378 -15712
rect -6866 -15752 -6378 -15746
rect -7158 -15820 -7148 -15796
rect -8132 -16352 -8126 -15822
rect -7154 -16350 -7148 -15820
rect -8132 -16372 -8118 -16352
rect -8902 -16422 -8414 -16416
rect -8902 -16456 -8890 -16422
rect -8426 -16456 -8414 -16422
rect -8902 -16462 -8414 -16456
rect -8692 -16524 -8632 -16462
rect -8902 -16530 -8414 -16524
rect -8902 -16564 -8890 -16530
rect -8426 -16564 -8414 -16530
rect -8902 -16570 -8414 -16564
rect -9198 -16646 -9184 -16614
rect -9190 -17168 -9184 -16646
rect -9198 -17190 -9184 -17168
rect -9150 -16646 -9138 -16614
rect -8178 -16614 -8118 -16372
rect -7158 -16372 -7148 -16350
rect -7114 -15820 -7098 -15796
rect -6140 -15796 -6080 -15554
rect -5120 -15554 -5112 -15526
rect -5078 -15004 -5060 -14978
rect -4108 -14978 -4048 -14736
rect -3086 -14736 -3076 -14722
rect -3042 -14184 -3026 -14160
rect -2066 -14160 -2006 -13918
rect -1050 -13918 -1040 -13890
rect -1006 -13366 -992 -13342
rect -30 -13342 30 -13100
rect -1006 -13890 -1000 -13366
rect -30 -13370 -22 -13342
rect -1006 -13918 -990 -13890
rect -1776 -13968 -1288 -13962
rect -1776 -14002 -1764 -13968
rect -1300 -14002 -1288 -13968
rect -1776 -14008 -1288 -14002
rect -1570 -14070 -1510 -14008
rect -1776 -14076 -1288 -14070
rect -1776 -14110 -1764 -14076
rect -1300 -14110 -1288 -14076
rect -1776 -14116 -1288 -14110
rect -2066 -14184 -2058 -14160
rect -3042 -14722 -3036 -14184
rect -2064 -14722 -2058 -14184
rect -3042 -14736 -3026 -14722
rect -3812 -14786 -3324 -14780
rect -3812 -14820 -3800 -14786
rect -3336 -14820 -3324 -14786
rect -3812 -14826 -3324 -14820
rect -3610 -14888 -3550 -14826
rect -3812 -14894 -3324 -14888
rect -3812 -14928 -3800 -14894
rect -3336 -14928 -3324 -14894
rect -3812 -14934 -3324 -14928
rect -5078 -15526 -5072 -15004
rect -4108 -15012 -4094 -14978
rect -5078 -15554 -5060 -15526
rect -4100 -15534 -4094 -15012
rect -5848 -15604 -5360 -15598
rect -5848 -15638 -5836 -15604
rect -5372 -15638 -5360 -15604
rect -5848 -15644 -5360 -15638
rect -5658 -15706 -5598 -15644
rect -5848 -15712 -5360 -15706
rect -5848 -15746 -5836 -15712
rect -5372 -15746 -5360 -15712
rect -5848 -15752 -5360 -15746
rect -7114 -16350 -7108 -15820
rect -6140 -15824 -6130 -15796
rect -7114 -16372 -7098 -16350
rect -6136 -16354 -6130 -15824
rect -7884 -16422 -7396 -16416
rect -7884 -16456 -7872 -16422
rect -7408 -16456 -7396 -16422
rect -7884 -16462 -7396 -16456
rect -7678 -16524 -7618 -16462
rect -7884 -16530 -7396 -16524
rect -7884 -16564 -7872 -16530
rect -7408 -16564 -7396 -16530
rect -7884 -16570 -7396 -16564
rect -8178 -16642 -8166 -16614
rect -9150 -17168 -9144 -16646
rect -8172 -17164 -8166 -16642
rect -9150 -17190 -9138 -17168
rect -9198 -17432 -9138 -17190
rect -8178 -17190 -8166 -17164
rect -8132 -16642 -8118 -16614
rect -7158 -16614 -7098 -16372
rect -6140 -16372 -6130 -16354
rect -6096 -15824 -6080 -15796
rect -5120 -15796 -5060 -15554
rect -4108 -15554 -4094 -15534
rect -4060 -15012 -4048 -14978
rect -3086 -14978 -3026 -14736
rect -2066 -14736 -2058 -14722
rect -2024 -14184 -2006 -14160
rect -1050 -14160 -990 -13918
rect -28 -13918 -22 -13370
rect 12 -13370 30 -13342
rect 12 -13894 18 -13370
rect 12 -13918 32 -13894
rect -758 -13968 -270 -13962
rect -758 -14002 -746 -13968
rect -282 -14002 -270 -13968
rect -758 -14008 -270 -14002
rect -550 -14070 -490 -14008
rect -758 -14076 -270 -14070
rect -758 -14110 -746 -14076
rect -282 -14110 -270 -14076
rect -758 -14116 -270 -14110
rect -1050 -14180 -1040 -14160
rect -2024 -14722 -2018 -14184
rect -1046 -14718 -1040 -14180
rect -2024 -14736 -2006 -14722
rect -2794 -14786 -2306 -14780
rect -2794 -14820 -2782 -14786
rect -2318 -14820 -2306 -14786
rect -2794 -14826 -2306 -14820
rect -2588 -14888 -2528 -14826
rect -2794 -14894 -2306 -14888
rect -2794 -14928 -2782 -14894
rect -2318 -14928 -2306 -14894
rect -2794 -14934 -2306 -14928
rect -3086 -15012 -3076 -14978
rect -4060 -15534 -4054 -15012
rect -3082 -15534 -3076 -15012
rect -4060 -15554 -4048 -15534
rect -4830 -15604 -4342 -15598
rect -4830 -15638 -4818 -15604
rect -4354 -15638 -4342 -15604
rect -4830 -15644 -4342 -15638
rect -4628 -15706 -4568 -15644
rect -4830 -15712 -4342 -15706
rect -4830 -15746 -4818 -15712
rect -4354 -15746 -4342 -15712
rect -4830 -15752 -4342 -15746
rect -5120 -15816 -5112 -15796
rect -6096 -16354 -6090 -15824
rect -5118 -16346 -5112 -15816
rect -6096 -16372 -6080 -16354
rect -6866 -16422 -6378 -16416
rect -6866 -16456 -6854 -16422
rect -6390 -16456 -6378 -16422
rect -6866 -16462 -6378 -16456
rect -6658 -16524 -6598 -16462
rect -6866 -16530 -6378 -16524
rect -6866 -16564 -6854 -16530
rect -6390 -16564 -6378 -16530
rect -6866 -16570 -6378 -16564
rect -7158 -16640 -7148 -16614
rect -8132 -17164 -8126 -16642
rect -7154 -17162 -7148 -16640
rect -8132 -17190 -8118 -17164
rect -8902 -17240 -8414 -17234
rect -8902 -17274 -8890 -17240
rect -8426 -17274 -8414 -17240
rect -8902 -17280 -8414 -17274
rect -8690 -17342 -8630 -17280
rect -8902 -17348 -8414 -17342
rect -8902 -17382 -8890 -17348
rect -8426 -17382 -8414 -17348
rect -8902 -17388 -8414 -17382
rect -9198 -17458 -9184 -17432
rect -9190 -17986 -9184 -17458
rect -9198 -18008 -9184 -17986
rect -9150 -17458 -9138 -17432
rect -8178 -17432 -8118 -17190
rect -7158 -17190 -7148 -17162
rect -7114 -16640 -7098 -16614
rect -6140 -16614 -6080 -16372
rect -5120 -16372 -5112 -16346
rect -5078 -15816 -5060 -15796
rect -4108 -15796 -4048 -15554
rect -3086 -15554 -3076 -15534
rect -3042 -15012 -3026 -14978
rect -2066 -14978 -2006 -14736
rect -1050 -14736 -1040 -14718
rect -1006 -14180 -990 -14160
rect -28 -14160 32 -13918
rect -1006 -14718 -1000 -14180
rect -1006 -14736 -990 -14718
rect -1776 -14786 -1288 -14780
rect -1776 -14820 -1764 -14786
rect -1300 -14820 -1288 -14786
rect -1776 -14826 -1288 -14820
rect -1576 -14888 -1516 -14826
rect -1776 -14894 -1288 -14888
rect -1776 -14928 -1764 -14894
rect -1300 -14928 -1288 -14894
rect -1776 -14934 -1288 -14928
rect -2066 -15012 -2058 -14978
rect -3042 -15534 -3036 -15012
rect -2064 -15534 -2058 -15012
rect -3042 -15554 -3026 -15534
rect -3812 -15604 -3324 -15598
rect -3812 -15638 -3800 -15604
rect -3336 -15638 -3324 -15604
rect -3812 -15644 -3324 -15638
rect -3612 -15706 -3552 -15644
rect -3812 -15712 -3324 -15706
rect -3812 -15746 -3800 -15712
rect -3336 -15746 -3324 -15712
rect -3812 -15752 -3324 -15746
rect -5078 -16346 -5072 -15816
rect -4108 -15824 -4094 -15796
rect -5078 -16372 -5060 -16346
rect -4100 -16354 -4094 -15824
rect -5848 -16422 -5360 -16416
rect -5848 -16456 -5836 -16422
rect -5372 -16456 -5360 -16422
rect -5848 -16462 -5360 -16456
rect -5656 -16524 -5596 -16462
rect -5848 -16530 -5360 -16524
rect -5848 -16564 -5836 -16530
rect -5372 -16564 -5360 -16530
rect -5848 -16570 -5360 -16564
rect -7114 -17162 -7108 -16640
rect -6140 -16644 -6130 -16614
rect -7114 -17190 -7098 -17162
rect -6136 -17166 -6130 -16644
rect -7884 -17240 -7396 -17234
rect -7884 -17274 -7872 -17240
rect -7408 -17274 -7396 -17240
rect -7884 -17280 -7396 -17274
rect -7676 -17342 -7616 -17280
rect -7884 -17348 -7396 -17342
rect -7884 -17382 -7872 -17348
rect -7408 -17382 -7396 -17348
rect -7884 -17388 -7396 -17382
rect -8178 -17454 -8166 -17432
rect -9150 -17986 -9144 -17458
rect -8172 -17982 -8166 -17454
rect -9150 -18008 -9138 -17986
rect -9198 -18250 -9138 -18008
rect -8178 -18008 -8166 -17982
rect -8132 -17454 -8118 -17432
rect -7158 -17432 -7098 -17190
rect -6140 -17190 -6130 -17166
rect -6096 -16644 -6080 -16614
rect -5120 -16614 -5060 -16372
rect -4108 -16372 -4094 -16354
rect -4060 -15824 -4048 -15796
rect -3086 -15796 -3026 -15554
rect -2066 -15554 -2058 -15534
rect -2024 -15012 -2006 -14978
rect -1050 -14978 -990 -14736
rect -28 -14736 -22 -14160
rect 12 -14184 32 -14160
rect 12 -14722 18 -14184
rect 12 -14736 32 -14722
rect -758 -14786 -270 -14780
rect -758 -14820 -746 -14786
rect -282 -14820 -270 -14786
rect -758 -14826 -270 -14820
rect -556 -14888 -496 -14826
rect -758 -14894 -270 -14888
rect -758 -14928 -746 -14894
rect -282 -14928 -270 -14894
rect -758 -14934 -270 -14928
rect -1050 -15008 -1040 -14978
rect -2024 -15534 -2018 -15012
rect -1046 -15530 -1040 -15008
rect -2024 -15554 -2006 -15534
rect -2794 -15604 -2306 -15598
rect -2794 -15638 -2782 -15604
rect -2318 -15638 -2306 -15604
rect -2794 -15644 -2306 -15638
rect -2590 -15706 -2530 -15644
rect -2794 -15712 -2306 -15706
rect -2794 -15746 -2782 -15712
rect -2318 -15746 -2306 -15712
rect -2794 -15752 -2306 -15746
rect -3086 -15824 -3076 -15796
rect -4060 -16354 -4054 -15824
rect -3082 -16354 -3076 -15824
rect -4060 -16372 -4048 -16354
rect -4830 -16422 -4342 -16416
rect -4830 -16456 -4818 -16422
rect -4354 -16456 -4342 -16422
rect -4830 -16462 -4342 -16456
rect -4626 -16524 -4566 -16462
rect -4830 -16530 -4342 -16524
rect -4830 -16564 -4818 -16530
rect -4354 -16564 -4342 -16530
rect -4830 -16570 -4342 -16564
rect -5120 -16636 -5112 -16614
rect -6096 -17166 -6090 -16644
rect -5118 -17158 -5112 -16636
rect -6096 -17190 -6080 -17166
rect -6866 -17240 -6378 -17234
rect -6866 -17274 -6854 -17240
rect -6390 -17274 -6378 -17240
rect -6866 -17280 -6378 -17274
rect -6656 -17342 -6596 -17280
rect -6866 -17348 -6378 -17342
rect -6866 -17382 -6854 -17348
rect -6390 -17382 -6378 -17348
rect -6866 -17388 -6378 -17382
rect -7158 -17452 -7148 -17432
rect -8132 -17982 -8126 -17454
rect -7154 -17980 -7148 -17452
rect -8132 -18008 -8118 -17982
rect -8902 -18058 -8414 -18052
rect -8902 -18092 -8890 -18058
rect -8426 -18092 -8414 -18058
rect -8902 -18098 -8414 -18092
rect -8688 -18160 -8628 -18098
rect -8902 -18166 -8414 -18160
rect -8902 -18200 -8890 -18166
rect -8426 -18200 -8414 -18166
rect -8902 -18206 -8414 -18200
rect -9198 -18276 -9184 -18250
rect -9190 -18826 -9184 -18276
rect -9150 -18276 -9138 -18250
rect -8178 -18250 -8118 -18008
rect -7158 -18008 -7148 -17980
rect -7114 -17452 -7098 -17432
rect -6140 -17432 -6080 -17190
rect -5120 -17190 -5112 -17158
rect -5078 -16636 -5060 -16614
rect -4108 -16614 -4048 -16372
rect -3086 -16372 -3076 -16354
rect -3042 -15824 -3026 -15796
rect -2066 -15796 -2006 -15554
rect -1050 -15554 -1040 -15530
rect -1006 -15008 -990 -14978
rect -28 -14978 32 -14736
rect -1006 -15530 -1000 -15008
rect -1006 -15554 -990 -15530
rect -1776 -15604 -1288 -15598
rect -1776 -15638 -1764 -15604
rect -1300 -15638 -1288 -15604
rect -1776 -15644 -1288 -15638
rect -1578 -15706 -1518 -15644
rect -1776 -15712 -1288 -15706
rect -1776 -15746 -1764 -15712
rect -1300 -15746 -1288 -15712
rect -1776 -15752 -1288 -15746
rect -2066 -15824 -2058 -15796
rect -3042 -16354 -3036 -15824
rect -2064 -16354 -2058 -15824
rect -3042 -16372 -3026 -16354
rect -3812 -16422 -3324 -16416
rect -3812 -16456 -3800 -16422
rect -3336 -16456 -3324 -16422
rect -3812 -16462 -3324 -16456
rect -3610 -16524 -3550 -16462
rect -3812 -16530 -3324 -16524
rect -3812 -16564 -3800 -16530
rect -3336 -16564 -3324 -16530
rect -3812 -16570 -3324 -16564
rect -5078 -17158 -5072 -16636
rect -4108 -16644 -4094 -16614
rect -5078 -17190 -5060 -17158
rect -4100 -17166 -4094 -16644
rect -5848 -17240 -5360 -17234
rect -5848 -17274 -5836 -17240
rect -5372 -17274 -5360 -17240
rect -5848 -17280 -5360 -17274
rect -5654 -17342 -5594 -17280
rect -5848 -17348 -5360 -17342
rect -5848 -17382 -5836 -17348
rect -5372 -17382 -5360 -17348
rect -5848 -17388 -5360 -17382
rect -7114 -17980 -7108 -17452
rect -6140 -17456 -6130 -17432
rect -7114 -18008 -7098 -17980
rect -6136 -17984 -6130 -17456
rect -7884 -18058 -7396 -18052
rect -7884 -18092 -7872 -18058
rect -7408 -18092 -7396 -18058
rect -7884 -18098 -7396 -18092
rect -7674 -18160 -7614 -18098
rect -7884 -18166 -7396 -18160
rect -7884 -18200 -7872 -18166
rect -7408 -18200 -7396 -18166
rect -7884 -18206 -7396 -18200
rect -8178 -18272 -8166 -18250
rect -9150 -18826 -9144 -18276
rect -9190 -18838 -9144 -18826
rect -8172 -18826 -8166 -18272
rect -8132 -18272 -8118 -18250
rect -7158 -18250 -7098 -18008
rect -6140 -18008 -6130 -17984
rect -6096 -17456 -6080 -17432
rect -5120 -17432 -5060 -17190
rect -4108 -17190 -4094 -17166
rect -4060 -16644 -4048 -16614
rect -3086 -16614 -3026 -16372
rect -2066 -16372 -2058 -16354
rect -2024 -15824 -2006 -15796
rect -1050 -15796 -990 -15554
rect -28 -15554 -22 -14978
rect 12 -15012 32 -14978
rect 12 -15534 18 -15012
rect 12 -15554 32 -15534
rect -758 -15604 -270 -15598
rect -758 -15638 -746 -15604
rect -282 -15638 -270 -15604
rect -758 -15644 -270 -15638
rect -558 -15706 -498 -15644
rect -758 -15712 -270 -15706
rect -758 -15746 -746 -15712
rect -282 -15746 -270 -15712
rect -758 -15752 -270 -15746
rect -1050 -15820 -1040 -15796
rect -2024 -16354 -2018 -15824
rect -1046 -16350 -1040 -15820
rect -2024 -16372 -2006 -16354
rect -2794 -16422 -2306 -16416
rect -2794 -16456 -2782 -16422
rect -2318 -16456 -2306 -16422
rect -2794 -16462 -2306 -16456
rect -2588 -16524 -2528 -16462
rect -2794 -16530 -2306 -16524
rect -2794 -16564 -2782 -16530
rect -2318 -16564 -2306 -16530
rect -2794 -16570 -2306 -16564
rect -3086 -16644 -3076 -16614
rect -4060 -17166 -4054 -16644
rect -3082 -17166 -3076 -16644
rect -4060 -17190 -4048 -17166
rect -4830 -17240 -4342 -17234
rect -4830 -17274 -4818 -17240
rect -4354 -17274 -4342 -17240
rect -4830 -17280 -4342 -17274
rect -4624 -17342 -4564 -17280
rect -4830 -17348 -4342 -17342
rect -4830 -17382 -4818 -17348
rect -4354 -17382 -4342 -17348
rect -4830 -17388 -4342 -17382
rect -5120 -17448 -5112 -17432
rect -6096 -17984 -6090 -17456
rect -5118 -17976 -5112 -17448
rect -6096 -18008 -6080 -17984
rect -6866 -18058 -6378 -18052
rect -6866 -18092 -6854 -18058
rect -6390 -18092 -6378 -18058
rect -6866 -18098 -6378 -18092
rect -6654 -18160 -6594 -18098
rect -6866 -18166 -6378 -18160
rect -6866 -18200 -6854 -18166
rect -6390 -18200 -6378 -18166
rect -6866 -18206 -6378 -18200
rect -7158 -18270 -7148 -18250
rect -8132 -18826 -8126 -18272
rect -7154 -18780 -7148 -18270
rect -8172 -18838 -8126 -18826
rect -7164 -18826 -7148 -18780
rect -7114 -18270 -7098 -18250
rect -6140 -18250 -6080 -18008
rect -5120 -18008 -5112 -17976
rect -5078 -17448 -5060 -17432
rect -4108 -17432 -4048 -17190
rect -3086 -17190 -3076 -17166
rect -3042 -16644 -3026 -16614
rect -2066 -16614 -2006 -16372
rect -1050 -16372 -1040 -16350
rect -1006 -15820 -990 -15796
rect -28 -15796 32 -15554
rect -1006 -16350 -1000 -15820
rect -1006 -16372 -990 -16350
rect -1776 -16422 -1288 -16416
rect -1776 -16456 -1764 -16422
rect -1300 -16456 -1288 -16422
rect -1776 -16462 -1288 -16456
rect -1576 -16524 -1516 -16462
rect -1776 -16530 -1288 -16524
rect -1776 -16564 -1764 -16530
rect -1300 -16564 -1288 -16530
rect -1776 -16570 -1288 -16564
rect -2066 -16644 -2058 -16614
rect -3042 -17166 -3036 -16644
rect -2064 -17166 -2058 -16644
rect -3042 -17190 -3026 -17166
rect -3812 -17240 -3324 -17234
rect -3812 -17274 -3800 -17240
rect -3336 -17274 -3324 -17240
rect -3812 -17280 -3324 -17274
rect -3608 -17342 -3548 -17280
rect -3812 -17348 -3324 -17342
rect -3812 -17382 -3800 -17348
rect -3336 -17382 -3324 -17348
rect -3812 -17388 -3324 -17382
rect -5078 -17976 -5072 -17448
rect -4108 -17456 -4094 -17432
rect -5078 -18008 -5060 -17976
rect -4100 -17984 -4094 -17456
rect -5848 -18058 -5360 -18052
rect -5848 -18092 -5836 -18058
rect -5372 -18092 -5360 -18058
rect -5848 -18098 -5360 -18092
rect -5652 -18160 -5592 -18098
rect -5848 -18166 -5360 -18160
rect -5848 -18200 -5836 -18166
rect -5372 -18200 -5360 -18166
rect -5848 -18206 -5360 -18200
rect -7114 -18780 -7108 -18270
rect -6140 -18274 -6130 -18250
rect -7114 -18826 -7104 -18780
rect -8902 -18876 -8414 -18870
rect -8902 -18910 -8890 -18876
rect -8426 -18910 -8414 -18876
rect -8902 -18916 -8414 -18910
rect -7884 -18876 -7396 -18870
rect -7884 -18910 -7872 -18876
rect -7408 -18910 -7396 -18876
rect -7884 -18916 -7672 -18910
rect -7612 -18916 -7396 -18910
rect -7164 -19000 -7104 -18826
rect -6136 -18826 -6130 -18274
rect -6096 -18274 -6080 -18250
rect -5120 -18250 -5060 -18008
rect -4108 -18008 -4094 -17984
rect -4060 -17456 -4048 -17432
rect -3086 -17432 -3026 -17190
rect -2066 -17190 -2058 -17166
rect -2024 -16644 -2006 -16614
rect -1050 -16614 -990 -16372
rect -28 -16372 -22 -15796
rect 12 -15824 32 -15796
rect 12 -16354 18 -15824
rect 12 -16372 32 -16354
rect -758 -16422 -270 -16416
rect -758 -16456 -746 -16422
rect -282 -16456 -270 -16422
rect -758 -16462 -270 -16456
rect -556 -16524 -496 -16462
rect -758 -16530 -270 -16524
rect -758 -16564 -746 -16530
rect -282 -16564 -270 -16530
rect -758 -16570 -270 -16564
rect -1050 -16640 -1040 -16614
rect -2024 -17166 -2018 -16644
rect -1046 -17162 -1040 -16640
rect -2024 -17190 -2006 -17166
rect -2794 -17240 -2306 -17234
rect -2794 -17274 -2782 -17240
rect -2318 -17274 -2306 -17240
rect -2794 -17280 -2306 -17274
rect -2586 -17342 -2526 -17280
rect -2794 -17348 -2306 -17342
rect -2794 -17382 -2782 -17348
rect -2318 -17382 -2306 -17348
rect -2794 -17388 -2306 -17382
rect -3086 -17456 -3076 -17432
rect -4060 -17984 -4054 -17456
rect -3082 -17984 -3076 -17456
rect -4060 -18008 -4048 -17984
rect -4830 -18058 -4342 -18052
rect -4830 -18092 -4818 -18058
rect -4354 -18092 -4342 -18058
rect -4830 -18098 -4342 -18092
rect -4622 -18160 -4562 -18098
rect -4830 -18166 -4342 -18160
rect -4830 -18200 -4818 -18166
rect -4354 -18200 -4342 -18166
rect -4830 -18206 -4342 -18200
rect -5120 -18266 -5112 -18250
rect -6096 -18826 -6090 -18274
rect -5118 -18778 -5112 -18266
rect -6136 -18838 -6090 -18826
rect -5126 -18826 -5112 -18778
rect -5078 -18266 -5060 -18250
rect -4108 -18250 -4048 -18008
rect -3086 -18008 -3076 -17984
rect -3042 -17456 -3026 -17432
rect -2066 -17432 -2006 -17190
rect -1050 -17190 -1040 -17162
rect -1006 -16640 -990 -16614
rect -28 -16614 32 -16372
rect -1006 -17162 -1000 -16640
rect -1006 -17190 -990 -17162
rect -1776 -17240 -1288 -17234
rect -1776 -17274 -1764 -17240
rect -1300 -17274 -1288 -17240
rect -1776 -17280 -1288 -17274
rect -1574 -17342 -1514 -17280
rect -1776 -17348 -1288 -17342
rect -1776 -17382 -1764 -17348
rect -1300 -17382 -1288 -17348
rect -1776 -17388 -1288 -17382
rect -2066 -17456 -2058 -17432
rect -3042 -17984 -3036 -17456
rect -2064 -17984 -2058 -17456
rect -3042 -18008 -3026 -17984
rect -3812 -18058 -3324 -18052
rect -3812 -18092 -3800 -18058
rect -3336 -18092 -3324 -18058
rect -3812 -18098 -3324 -18092
rect -3606 -18160 -3546 -18098
rect -3812 -18166 -3324 -18160
rect -3812 -18200 -3800 -18166
rect -3336 -18200 -3324 -18166
rect -3812 -18206 -3324 -18200
rect -5078 -18778 -5072 -18266
rect -4108 -18274 -4094 -18250
rect -5078 -18826 -5066 -18778
rect -6866 -18876 -6378 -18870
rect -6866 -18910 -6854 -18876
rect -6390 -18910 -6378 -18876
rect -6866 -18916 -6378 -18910
rect -5848 -18876 -5360 -18870
rect -5848 -18910 -5836 -18876
rect -5372 -18910 -5360 -18876
rect -5848 -18916 -5360 -18910
rect -5126 -19000 -5066 -18826
rect -4100 -18826 -4094 -18274
rect -4060 -18274 -4048 -18250
rect -3086 -18250 -3026 -18008
rect -2066 -18008 -2058 -17984
rect -2024 -17456 -2006 -17432
rect -1050 -17432 -990 -17190
rect -28 -17190 -22 -16614
rect 12 -16644 32 -16614
rect 12 -17166 18 -16644
rect 12 -17190 32 -17166
rect -758 -17240 -270 -17234
rect -758 -17274 -746 -17240
rect -282 -17274 -270 -17240
rect -758 -17280 -270 -17274
rect -554 -17342 -494 -17280
rect -758 -17348 -270 -17342
rect -758 -17382 -746 -17348
rect -282 -17382 -270 -17348
rect -758 -17388 -270 -17382
rect -1050 -17452 -1040 -17432
rect -2024 -17984 -2018 -17456
rect -1046 -17980 -1040 -17452
rect -2024 -18008 -2006 -17984
rect -2794 -18058 -2306 -18052
rect -2794 -18092 -2782 -18058
rect -2318 -18092 -2306 -18058
rect -2794 -18098 -2306 -18092
rect -2584 -18160 -2524 -18098
rect -2794 -18166 -2306 -18160
rect -2794 -18200 -2782 -18166
rect -2318 -18200 -2306 -18166
rect -2794 -18206 -2306 -18200
rect -3086 -18274 -3076 -18250
rect -4060 -18826 -4054 -18274
rect -3082 -18782 -3076 -18274
rect -4100 -18838 -4054 -18826
rect -3090 -18826 -3076 -18782
rect -3042 -18274 -3026 -18250
rect -2066 -18250 -2006 -18008
rect -1050 -18008 -1040 -17980
rect -1006 -17452 -990 -17432
rect -28 -17432 32 -17190
rect -1006 -17980 -1000 -17452
rect -1006 -18008 -990 -17980
rect -1776 -18058 -1288 -18052
rect -1776 -18092 -1764 -18058
rect -1300 -18092 -1288 -18058
rect -1776 -18098 -1288 -18092
rect -1572 -18160 -1512 -18098
rect -1776 -18166 -1288 -18160
rect -1776 -18200 -1764 -18166
rect -1300 -18200 -1288 -18166
rect -1776 -18206 -1288 -18200
rect -2066 -18274 -2058 -18250
rect -3042 -18782 -3036 -18274
rect -3042 -18826 -3030 -18782
rect -4830 -18876 -4342 -18870
rect -4830 -18910 -4818 -18876
rect -4354 -18910 -4342 -18876
rect -4830 -18916 -4342 -18910
rect -3812 -18876 -3324 -18870
rect -3812 -18910 -3800 -18876
rect -3336 -18910 -3324 -18876
rect -3812 -18916 -3324 -18910
rect -3090 -19000 -3030 -18826
rect -2064 -18826 -2058 -18274
rect -2024 -18274 -2006 -18250
rect -1050 -18250 -990 -18008
rect -28 -18008 -22 -17432
rect 12 -17456 32 -17432
rect 12 -17984 18 -17456
rect 12 -18008 32 -17984
rect -758 -18058 -270 -18052
rect -758 -18092 -746 -18058
rect -282 -18092 -270 -18058
rect -758 -18098 -270 -18092
rect -552 -18160 -492 -18098
rect -758 -18166 -270 -18160
rect -758 -18200 -746 -18166
rect -282 -18200 -270 -18166
rect -758 -18206 -270 -18200
rect -1050 -18270 -1040 -18250
rect -2024 -18826 -2018 -18274
rect -1046 -18784 -1040 -18270
rect -2064 -18838 -2018 -18826
rect -1054 -18826 -1040 -18784
rect -1006 -18270 -990 -18250
rect -28 -18250 32 -18008
rect -1006 -18784 -1000 -18270
rect -28 -18772 -22 -18250
rect -1006 -18826 -994 -18784
rect -2794 -18876 -2306 -18870
rect -2794 -18910 -2782 -18876
rect -2318 -18910 -2306 -18876
rect -2794 -18916 -2306 -18910
rect -1776 -18876 -1288 -18870
rect -1776 -18910 -1764 -18876
rect -1300 -18910 -1288 -18876
rect -1776 -18916 -1288 -18910
rect -1054 -19000 -994 -18826
rect -34 -18826 -22 -18772
rect 12 -18274 32 -18250
rect 12 -18772 18 -18274
rect 12 -18826 26 -18772
rect 1150 -18822 1210 -11682
rect -758 -18876 -270 -18870
rect -758 -18910 -746 -18876
rect -282 -18910 -270 -18876
rect -758 -18916 -270 -18910
rect -540 -19000 -480 -18916
rect -34 -19000 26 -18826
rect 1144 -18882 1150 -18822
rect 1210 -18882 1216 -18822
rect -7164 -19060 1130 -19000
rect -3404 -19808 -3398 -19748
rect -3338 -19808 -3332 -19748
rect -9508 -19894 -9448 -19888
rect -5434 -19954 -5428 -19894
rect -5368 -19954 -5362 -19894
rect -10668 -20082 -10662 -20022
rect -10602 -20082 -10596 -20022
rect -10662 -22254 -10602 -20082
rect -9508 -20086 -9448 -19954
rect -7990 -20082 -7984 -20022
rect -7924 -20082 -7918 -20022
rect -6958 -20082 -6952 -20022
rect -6892 -20082 -6886 -20022
rect -10524 -20146 -9448 -20086
rect -10524 -20320 -10464 -20146
rect -10016 -20228 -9956 -20146
rect -9508 -20314 -9448 -20146
rect -7984 -20224 -7924 -20082
rect -6952 -20220 -6892 -20082
rect -5428 -20338 -5368 -19954
rect -3898 -20082 -3892 -20022
rect -3832 -20082 -3826 -20022
rect -3892 -20220 -3832 -20082
rect -9004 -20984 -8944 -20904
rect -9010 -21044 -9004 -20984
rect -8944 -21044 -8938 -20984
rect -9510 -21148 -9504 -21088
rect -9444 -21148 -9438 -21088
rect -9504 -21190 -9444 -21148
rect -10524 -21250 -9444 -21190
rect -10524 -21432 -10464 -21250
rect -10020 -21328 -9960 -21250
rect -10668 -22314 -10662 -22254
rect -10602 -22314 -10596 -22254
rect -10662 -24380 -10602 -22314
rect -9504 -22570 -9444 -21250
rect -8486 -21192 -8426 -20786
rect -7986 -21044 -7980 -20984
rect -7920 -21044 -7914 -20984
rect -9012 -22254 -8952 -22010
rect -9018 -22314 -9012 -22254
rect -8952 -22314 -8946 -22254
rect -9012 -22450 -8952 -22314
rect -10520 -23206 -10460 -23040
rect -10028 -23206 -9968 -23120
rect -9500 -23206 -9440 -23044
rect -10520 -23266 -9440 -23206
rect -9500 -23306 -9440 -23266
rect -8486 -23198 -8426 -21252
rect -7980 -21340 -7920 -21044
rect -7468 -21088 -7408 -20804
rect -6954 -21044 -6948 -20984
rect -6888 -21044 -6882 -20984
rect -7474 -21148 -7468 -21088
rect -7408 -21148 -7402 -21088
rect -6948 -21336 -6888 -21044
rect -6450 -21192 -6390 -20788
rect -5948 -20984 -5888 -20902
rect -4928 -20984 -4868 -20902
rect -5954 -21044 -5948 -20984
rect -5888 -21044 -5882 -20984
rect -4934 -21044 -4928 -20984
rect -4868 -21044 -4862 -20984
rect -5438 -21148 -5432 -21088
rect -5372 -21148 -5366 -21088
rect -7474 -22134 -7414 -21924
rect -7480 -22194 -7474 -22134
rect -7414 -22194 -7408 -22134
rect -7474 -22568 -7414 -22194
rect -9506 -23366 -9500 -23306
rect -9440 -23366 -9434 -23306
rect -9012 -23478 -9006 -23418
rect -8946 -23478 -8940 -23418
rect -9006 -23558 -8946 -23478
rect -8486 -23712 -8426 -23258
rect -7982 -23418 -7922 -23122
rect -7470 -23366 -7464 -23306
rect -7404 -23366 -7398 -23306
rect -7988 -23478 -7982 -23418
rect -7922 -23478 -7916 -23418
rect -7464 -23650 -7404 -23366
rect -6950 -23418 -6890 -23126
rect -6450 -23198 -6390 -21252
rect -5942 -22254 -5882 -22012
rect -5948 -22314 -5942 -22254
rect -5882 -22314 -5876 -22254
rect -5942 -22448 -5882 -22314
rect -5432 -22604 -5372 -21148
rect -4418 -21192 -4358 -20778
rect -3914 -21044 -3908 -20984
rect -3848 -21044 -3842 -20984
rect -4424 -21252 -4418 -21192
rect -4358 -21252 -4352 -21192
rect -4934 -22254 -4874 -22010
rect -4940 -22314 -4934 -22254
rect -4874 -22314 -4868 -22254
rect -4934 -22448 -4874 -22314
rect -6956 -23478 -6950 -23418
rect -6890 -23478 -6884 -23418
rect -6450 -23648 -6390 -23258
rect -5428 -23306 -5368 -23012
rect -4418 -23198 -4358 -21252
rect -3908 -21330 -3848 -21044
rect -3398 -21088 -3338 -19808
rect -1374 -19954 -1368 -19894
rect -1308 -19954 -1302 -19894
rect 810 -19954 816 -19894
rect 876 -19954 882 -19894
rect -2902 -20082 -2896 -20022
rect -2836 -20082 -2830 -20022
rect -2896 -20232 -2836 -20082
rect -1368 -20306 -1308 -19954
rect -2898 -20984 -2838 -20978
rect -3404 -21148 -3398 -21088
rect -3338 -21148 -3332 -21088
rect -2898 -21340 -2838 -21044
rect -2384 -21192 -2324 -20788
rect -1884 -20984 -1824 -20900
rect -866 -20984 -806 -20902
rect -1890 -21044 -1884 -20984
rect -1824 -21044 -1818 -20984
rect -866 -21050 -806 -21044
rect -340 -21078 -280 -20816
rect 164 -21078 224 -20896
rect 676 -21078 736 -20796
rect -1368 -21148 -1362 -21088
rect -1302 -21148 -1296 -21088
rect -340 -21138 736 -21078
rect -3398 -22134 -3338 -21906
rect -3404 -22194 -3398 -22134
rect -3338 -22194 -3332 -22134
rect -3398 -22540 -3338 -22194
rect -5434 -23366 -5428 -23306
rect -5368 -23366 -5362 -23306
rect -5956 -23478 -5950 -23418
rect -5890 -23478 -5884 -23418
rect -4936 -23478 -4930 -23418
rect -4870 -23478 -4864 -23418
rect -5950 -23560 -5890 -23478
rect -4930 -23560 -4870 -23478
rect -4418 -23670 -4358 -23258
rect -3910 -23418 -3850 -23132
rect -3400 -23366 -3394 -23306
rect -3334 -23366 -3328 -23306
rect -3916 -23478 -3910 -23418
rect -3850 -23478 -3844 -23418
rect -3394 -23656 -3334 -23366
rect -2900 -23418 -2840 -23122
rect -2900 -23484 -2840 -23478
rect -2384 -23198 -2324 -21252
rect -1872 -22254 -1812 -22018
rect -1878 -22314 -1872 -22254
rect -1812 -22314 -1806 -22254
rect -1872 -22444 -1812 -22314
rect -1362 -22554 -1302 -21148
rect -340 -21192 -280 -21138
rect -846 -22254 -786 -22010
rect -340 -22198 -280 -21252
rect 164 -21332 224 -21138
rect 160 -22198 220 -22012
rect 676 -22198 736 -21138
rect 816 -22134 876 -19954
rect 930 -21044 936 -20984
rect 996 -21044 1002 -20984
rect 810 -22194 816 -22134
rect 876 -22194 882 -22134
rect -852 -22314 -846 -22254
rect -786 -22314 -780 -22254
rect -340 -22258 736 -22198
rect -846 -22450 -786 -22314
rect -2384 -23652 -2324 -23258
rect -1358 -23306 -1298 -23028
rect -340 -23198 -280 -22258
rect 160 -22452 220 -22258
rect -346 -23258 -340 -23198
rect -280 -23258 -274 -23198
rect -1364 -23366 -1358 -23306
rect -1298 -23366 -1292 -23306
rect -340 -23310 -280 -23258
rect 168 -23310 228 -23120
rect 676 -23310 736 -22258
rect -340 -23370 736 -23310
rect -868 -23418 -808 -23412
rect -1892 -23478 -1886 -23418
rect -1826 -23478 -1820 -23418
rect -1886 -23562 -1826 -23478
rect -868 -23560 -808 -23478
rect -340 -23674 -280 -23370
rect 168 -23560 228 -23370
rect 676 -23652 736 -23370
rect -10524 -24330 -10464 -24144
rect -10020 -24330 -9960 -24244
rect -9506 -24330 -9446 -24150
rect -10668 -24440 -10662 -24380
rect -10602 -24440 -10596 -24380
rect -10524 -24390 -9446 -24330
rect -7992 -24380 -7932 -24238
rect -6960 -24380 -6900 -24242
rect -9506 -24510 -9446 -24390
rect -7998 -24440 -7992 -24380
rect -7932 -24440 -7926 -24380
rect -6966 -24440 -6960 -24380
rect -6900 -24440 -6894 -24380
rect -5426 -24510 -5366 -24126
rect -3900 -24380 -3840 -24242
rect -2904 -24380 -2844 -24230
rect -3906 -24440 -3900 -24380
rect -3840 -24440 -3834 -24380
rect -2910 -24440 -2904 -24380
rect -2844 -24440 -2838 -24380
rect -1366 -24510 -1306 -24158
rect 816 -24510 876 -22194
rect 936 -23418 996 -21044
rect 930 -23478 936 -23418
rect 996 -23478 1002 -23418
rect -5432 -24570 -5426 -24510
rect -5366 -24570 -5360 -24510
rect -1372 -24570 -1366 -24510
rect -1306 -24570 -1300 -24510
rect 810 -24570 816 -24510
rect 876 -24570 882 -24510
rect -9506 -24576 -9446 -24570
rect -10064 -24976 172 -24916
rect -10064 -25186 -10004 -24976
rect -9564 -25098 -9504 -24976
rect -9042 -25196 -8982 -24976
rect -8544 -25098 -8484 -24976
rect -7510 -25104 -7450 -24976
rect -6488 -25104 -6428 -24976
rect -5498 -25104 -5438 -24976
rect -4974 -25194 -4914 -24976
rect -4464 -25110 -4404 -24976
rect -3474 -25098 -3414 -24976
rect -2442 -25110 -2382 -24976
rect -1438 -25098 -1378 -24976
rect -898 -25220 -838 -24976
rect -418 -25104 -358 -24976
rect 112 -25192 172 -24976
rect -8028 -25876 -7968 -25670
rect -8034 -25936 -8028 -25876
rect -7968 -25936 -7962 -25876
rect -12328 -27116 -12216 -26330
rect -8028 -26430 -7968 -25936
rect -7010 -25988 -6950 -25694
rect -5990 -25876 -5930 -25682
rect -3954 -25876 -3894 -25682
rect -5996 -25936 -5990 -25876
rect -5930 -25936 -5924 -25876
rect -3960 -25936 -3954 -25876
rect -3894 -25936 -3888 -25876
rect -7016 -26048 -7010 -25988
rect -6950 -26048 -6944 -25988
rect -5990 -26430 -5930 -25936
rect -3954 -26430 -3894 -25936
rect -2936 -25988 -2876 -25690
rect -1918 -25876 -1858 -25696
rect -1924 -25936 -1918 -25876
rect -1858 -25936 -1852 -25876
rect -2942 -26048 -2936 -25988
rect -2876 -26048 -2870 -25988
rect -1918 -26430 -1858 -25936
rect 1070 -25988 1130 -19060
rect 1282 -19894 1342 -11554
rect 1276 -19954 1282 -19894
rect 1342 -19954 1348 -19894
rect 1402 -20022 1462 -11552
rect 1396 -20082 1402 -20022
rect 1462 -20082 1468 -20022
rect 1542 -20984 1602 -11534
rect 1654 -11672 1660 -11612
rect 1720 -11672 1726 -11612
rect 1660 -17740 1720 -11672
rect 1770 -12354 1830 -11518
rect 1764 -12414 1770 -12354
rect 1830 -12414 1836 -12354
rect 1888 -15274 1948 -11418
rect 2216 -12220 2276 -11408
rect 2210 -12280 2216 -12220
rect 2276 -12280 2282 -12220
rect 2006 -13638 2012 -13578
rect 2072 -13638 2078 -13578
rect 1886 -15280 1948 -15274
rect 1946 -15340 1948 -15280
rect 1886 -15346 1948 -15340
rect 1654 -17800 1660 -17740
rect 1720 -17800 1726 -17740
rect 1536 -21044 1542 -20984
rect 1602 -21044 1608 -20984
rect 1888 -21342 1948 -15346
rect 2012 -16274 2072 -13638
rect 2218 -13974 2224 -13914
rect 2284 -13974 2290 -13914
rect 2114 -15234 2120 -15174
rect 2180 -15234 2186 -15174
rect 2006 -16334 2012 -16274
rect 2072 -16334 2078 -16274
rect 2120 -21192 2180 -15234
rect 2224 -16510 2284 -13974
rect 2336 -16396 2396 -11416
rect 2442 -11492 2502 -11486
rect 2442 -14036 2502 -11552
rect 13248 -11848 13254 -11842
rect 2568 -11902 13254 -11848
rect 13314 -11848 13320 -11842
rect 18352 -11848 18358 -11842
rect 13314 -11902 18358 -11848
rect 18418 -11848 18424 -11842
rect 22418 -11848 22478 -11842
rect 18418 -11902 22418 -11848
rect 2568 -11908 22418 -11902
rect 22478 -11908 22990 -11848
rect 2568 -13914 2628 -11908
rect 3090 -11996 3150 -11908
rect 4100 -12010 4160 -11908
rect 3080 -12828 3140 -12672
rect 3586 -13578 3646 -12590
rect 4086 -12822 4146 -12666
rect 4606 -12924 4666 -11908
rect 5130 -11992 5190 -11908
rect 6142 -12010 6202 -11908
rect 5098 -12816 5158 -12660
rect 5620 -13580 5680 -12578
rect 6120 -12828 6180 -12672
rect 6638 -12928 6698 -11908
rect 7154 -11992 7214 -11908
rect 8154 -11998 8214 -11908
rect 7132 -12828 7192 -12672
rect 7656 -13580 7716 -12584
rect 8162 -12828 8222 -12672
rect 8676 -12908 8736 -11908
rect 9188 -12004 9248 -11908
rect 10200 -12004 10260 -11908
rect 9168 -12822 9228 -12666
rect 9694 -13580 9754 -12584
rect 10190 -12822 10250 -12666
rect 10712 -12916 10772 -11908
rect 11224 -12004 11284 -11908
rect 12236 -11992 12296 -11908
rect 11214 -12828 11274 -12672
rect 11732 -13580 11792 -12578
rect 12220 -12822 12280 -12666
rect 12744 -12914 12804 -11908
rect 13258 -11998 13318 -11908
rect 14270 -12010 14330 -11908
rect 13244 -12816 13304 -12660
rect 13766 -13580 13826 -12578
rect 14266 -12822 14326 -12666
rect 14782 -12916 14842 -11908
rect 15294 -12010 15354 -11908
rect 16312 -11998 16372 -11908
rect 15278 -12822 15338 -12666
rect 15802 -13580 15862 -12578
rect 16290 -12828 16350 -12672
rect 16818 -12890 16878 -11908
rect 17334 -11992 17394 -11908
rect 18358 -11992 18418 -11908
rect 17314 -12816 17374 -12660
rect 17840 -13580 17900 -12554
rect 18336 -12834 18396 -12678
rect 18854 -12908 18914 -11908
rect 19376 -11998 19436 -11908
rect 20388 -11998 20448 -11908
rect 19354 -12822 19414 -12666
rect 19874 -13580 19934 -12514
rect 20384 -12810 20444 -12654
rect 20892 -12908 20952 -11908
rect 21398 -11992 21458 -11908
rect 22416 -11914 22478 -11908
rect 22416 -12004 22476 -11914
rect 21396 -12810 21456 -12654
rect 21910 -13580 21970 -12564
rect 22396 -12828 22456 -12672
rect 22930 -12716 22990 -11908
rect 24816 -12070 24928 -11284
rect 22930 -12776 23710 -12716
rect 22930 -12916 22990 -12776
rect 3646 -13638 23588 -13580
rect 3586 -13640 23588 -13638
rect 3586 -13644 3646 -13640
rect 4594 -13854 4600 -13794
rect 4660 -13854 4666 -13794
rect 6634 -13854 6640 -13794
rect 6700 -13854 6706 -13794
rect 8674 -13854 8680 -13794
rect 8740 -13854 8746 -13794
rect 10704 -13854 10710 -13794
rect 10770 -13854 10776 -13794
rect 12744 -13854 12750 -13794
rect 12810 -13854 12816 -13794
rect 14776 -13854 14782 -13794
rect 14842 -13854 14848 -13794
rect 16816 -13854 16822 -13794
rect 16882 -13854 16888 -13794
rect 18852 -13854 18858 -13794
rect 18918 -13854 18924 -13794
rect 20886 -13854 20892 -13794
rect 20952 -13854 20958 -13794
rect 2562 -13974 2568 -13914
rect 2628 -13974 2634 -13914
rect 4086 -13980 4092 -13920
rect 4152 -13980 4158 -13920
rect 2436 -14096 2442 -14036
rect 2502 -14096 2508 -14036
rect 2442 -16170 2502 -14096
rect 2864 -14160 3076 -14154
rect 3136 -14160 3352 -14154
rect 4092 -14160 4152 -13980
rect 2864 -14194 2876 -14160
rect 3340 -14194 3352 -14160
rect 2864 -14200 3352 -14194
rect 4600 -14244 4660 -13854
rect 5106 -13920 5166 -13914
rect 5106 -14160 5166 -13980
rect 6128 -13920 6188 -13914
rect 6128 -14160 6188 -13980
rect 5630 -14244 5676 -14232
rect 2568 -14278 2582 -14244
rect 2576 -14770 2582 -14278
rect 2568 -14820 2582 -14770
rect 2616 -14278 2628 -14244
rect 2616 -14770 2622 -14278
rect 3586 -14292 3600 -14244
rect 2616 -14820 2628 -14770
rect 3594 -14784 3600 -14292
rect 2568 -14958 2628 -14820
rect 3586 -14820 3600 -14784
rect 3634 -14292 3646 -14244
rect 3634 -14784 3640 -14292
rect 4600 -14312 4618 -14244
rect 4612 -14756 4618 -14312
rect 3634 -14820 3646 -14784
rect 2864 -14870 3352 -14864
rect 2864 -14904 2876 -14870
rect 3340 -14904 3352 -14870
rect 2864 -14910 3352 -14904
rect 3070 -14958 3130 -14910
rect 3586 -14958 3646 -14820
rect 4604 -14820 4618 -14756
rect 4652 -14276 4664 -14244
rect 4652 -14312 4660 -14276
rect 4652 -14756 4658 -14312
rect 4652 -14820 4664 -14756
rect 5630 -14774 5636 -14244
rect 5626 -14792 5636 -14774
rect 5624 -14820 5636 -14792
rect 5670 -14774 5676 -14244
rect 6640 -14244 6700 -13854
rect 7142 -13920 7202 -13914
rect 7140 -13980 7142 -13974
rect 8168 -13920 8228 -13914
rect 7140 -13986 7202 -13980
rect 8166 -13980 8168 -13974
rect 8166 -13986 8228 -13980
rect 7140 -14160 7200 -13986
rect 7650 -14096 7656 -14036
rect 7716 -14096 7722 -14036
rect 6640 -14298 6654 -14244
rect 6648 -14748 6654 -14298
rect 6644 -14772 6654 -14748
rect 5670 -14820 5686 -14774
rect 6642 -14820 6654 -14772
rect 6688 -14298 6700 -14244
rect 7656 -14244 7716 -14096
rect 8166 -14160 8226 -13986
rect 7656 -14286 7672 -14244
rect 6688 -14748 6694 -14298
rect 7666 -14744 7672 -14286
rect 6688 -14820 6704 -14748
rect 7656 -14820 7672 -14744
rect 7706 -14286 7716 -14244
rect 8680 -14244 8740 -13854
rect 9180 -13920 9240 -13914
rect 9180 -14160 9240 -13980
rect 10216 -13920 10276 -13914
rect 10216 -14160 10276 -13980
rect 10710 -14244 10770 -13854
rect 11222 -13920 11282 -13914
rect 12230 -13980 12236 -13920
rect 12296 -13980 12302 -13920
rect 11222 -14160 11282 -13980
rect 12236 -14160 12296 -13980
rect 12750 -14244 12810 -13854
rect 13252 -13920 13312 -13914
rect 13252 -14160 13312 -13980
rect 14260 -13920 14320 -13914
rect 14320 -13980 14322 -13974
rect 14260 -13986 14322 -13980
rect 14262 -14160 14322 -13986
rect 14782 -14244 14842 -13854
rect 15276 -13920 15336 -13914
rect 16300 -13920 16360 -13914
rect 15336 -13980 15338 -13974
rect 15276 -13986 15338 -13980
rect 15278 -14160 15338 -13986
rect 16300 -14160 16360 -13980
rect 16822 -14244 16882 -13854
rect 17322 -13920 17382 -13914
rect 18344 -13920 18404 -13914
rect 17322 -14160 17382 -13980
rect 18342 -13980 18344 -13974
rect 18342 -13986 18404 -13980
rect 17838 -14096 17844 -14036
rect 17904 -14096 17910 -14036
rect 7706 -14744 7712 -14286
rect 8680 -14318 8690 -14244
rect 7706 -14760 7716 -14744
rect 7706 -14820 7720 -14760
rect 8684 -14764 8690 -14318
rect 8676 -14820 8690 -14764
rect 8724 -14318 8740 -14244
rect 9696 -14294 9708 -14244
rect 8724 -14764 8730 -14318
rect 9702 -14756 9708 -14294
rect 8724 -14820 8736 -14764
rect 9696 -14784 9708 -14756
rect 9694 -14820 9708 -14784
rect 9742 -14294 9756 -14244
rect 9742 -14756 9748 -14294
rect 10710 -14312 10726 -14244
rect 10720 -14744 10726 -14312
rect 9742 -14820 9756 -14756
rect 3882 -14870 4370 -14864
rect 3882 -14904 3894 -14870
rect 4358 -14904 4370 -14870
rect 3882 -14910 4370 -14904
rect 2568 -15018 3646 -14958
rect 3586 -15174 3646 -15018
rect 4096 -15068 4156 -14910
rect 4604 -14958 4664 -14820
rect 4900 -14870 5388 -14864
rect 4900 -14904 4912 -14870
rect 5376 -14904 5388 -14870
rect 4900 -14910 5388 -14904
rect 4598 -15018 4604 -14958
rect 4664 -15018 4670 -14958
rect 4090 -15128 4096 -15068
rect 4156 -15128 4162 -15068
rect 3580 -15234 3586 -15174
rect 3646 -15234 3652 -15174
rect 2566 -15340 2572 -15280
rect 2632 -15340 2638 -15280
rect 3064 -15340 3070 -15280
rect 3130 -15340 3136 -15280
rect 3576 -15340 3582 -15280
rect 3642 -15340 3648 -15280
rect 2572 -15476 2632 -15340
rect 3070 -15386 3130 -15340
rect 2864 -15392 3352 -15386
rect 2864 -15426 2876 -15392
rect 3340 -15426 3352 -15392
rect 2864 -15432 3352 -15426
rect 2572 -15516 2582 -15476
rect 2576 -16052 2582 -15516
rect 2616 -15516 2632 -15476
rect 3582 -15476 3642 -15340
rect 4096 -15386 4156 -15128
rect 3882 -15392 4370 -15386
rect 3882 -15426 3894 -15392
rect 4358 -15426 4370 -15392
rect 3882 -15432 4370 -15426
rect 2616 -16052 2622 -15516
rect 3582 -15522 3600 -15476
rect 2576 -16064 2622 -16052
rect 3594 -16052 3600 -15522
rect 3634 -15522 3642 -15476
rect 4604 -15476 4664 -15018
rect 5118 -15068 5178 -14910
rect 5112 -15128 5118 -15068
rect 5178 -15128 5184 -15068
rect 5118 -15386 5178 -15128
rect 5626 -15174 5686 -14820
rect 5918 -14870 6406 -14864
rect 5918 -14904 5930 -14870
rect 6394 -14904 6406 -14870
rect 5918 -14910 6272 -14904
rect 6332 -14910 6406 -14904
rect 6132 -15068 6192 -14910
rect 6644 -14958 6704 -14820
rect 6936 -14870 7424 -14864
rect 6936 -14904 6948 -14870
rect 7412 -14904 7424 -14870
rect 6936 -14910 7144 -14904
rect 7146 -14910 7424 -14904
rect 7954 -14870 8442 -14864
rect 7954 -14904 7966 -14870
rect 8430 -14904 8442 -14870
rect 7954 -14910 8224 -14904
rect 8244 -14910 8442 -14904
rect 6638 -15018 6644 -14958
rect 6704 -15018 6710 -14958
rect 6126 -15128 6132 -15068
rect 6192 -15128 6198 -15068
rect 5620 -15234 5626 -15174
rect 5686 -15234 5692 -15174
rect 6132 -15386 6192 -15128
rect 4900 -15392 5388 -15386
rect 4900 -15426 4912 -15392
rect 5376 -15426 5388 -15392
rect 4900 -15432 5388 -15426
rect 5918 -15392 6192 -15386
rect 6196 -15392 6406 -15386
rect 5918 -15426 5930 -15392
rect 6394 -15426 6406 -15392
rect 5918 -15432 6406 -15426
rect 6644 -15476 6704 -15018
rect 7146 -15068 7206 -14910
rect 8164 -15068 8224 -14910
rect 8676 -14958 8736 -14820
rect 8972 -14870 9460 -14864
rect 8972 -14904 8984 -14870
rect 9448 -14904 9460 -14870
rect 8972 -14910 9460 -14904
rect 8670 -15018 8676 -14958
rect 8736 -15018 8742 -14958
rect 7140 -15128 7146 -15068
rect 7206 -15128 7212 -15068
rect 8158 -15128 8164 -15068
rect 8224 -15128 8230 -15068
rect 7146 -15386 7206 -15128
rect 7650 -15234 7656 -15174
rect 7716 -15234 7722 -15174
rect 6936 -15392 7138 -15386
rect 7146 -15392 7424 -15386
rect 6936 -15426 6948 -15392
rect 7412 -15426 7424 -15392
rect 6936 -15432 7424 -15426
rect 4604 -15514 4618 -15476
rect 3634 -16052 3640 -15522
rect 4612 -15994 4618 -15514
rect 3594 -16064 3640 -16052
rect 4598 -16052 4618 -15994
rect 4652 -15514 4664 -15476
rect 4652 -16052 4658 -15514
rect 5624 -15528 5636 -15476
rect 5630 -16032 5636 -15528
rect 2864 -16102 3352 -16096
rect 2864 -16136 2876 -16102
rect 3340 -16136 3352 -16102
rect 2864 -16142 3352 -16136
rect 3882 -16102 4370 -16096
rect 3882 -16136 3894 -16102
rect 4358 -16136 4370 -16102
rect 3882 -16142 4370 -16136
rect 2436 -16230 2442 -16170
rect 2502 -16230 2508 -16170
rect 4598 -16274 4658 -16052
rect 5620 -16052 5636 -16032
rect 5670 -15528 5684 -15476
rect 5670 -16032 5676 -15528
rect 6642 -15540 6654 -15476
rect 6648 -15988 6654 -15540
rect 5670 -16052 5680 -16032
rect 4900 -16102 5388 -16096
rect 4900 -16136 4912 -16102
rect 5376 -16136 5388 -16102
rect 4900 -16142 5388 -16136
rect 2560 -16334 2566 -16274
rect 2626 -16334 2632 -16274
rect 4080 -16334 4086 -16274
rect 4146 -16334 4152 -16274
rect 4592 -16334 4598 -16274
rect 4658 -16334 4664 -16274
rect 2330 -16456 2336 -16396
rect 2396 -16456 2402 -16396
rect 2218 -16570 2224 -16510
rect 2284 -16570 2290 -16510
rect 2336 -17638 2396 -16456
rect 2566 -16710 2626 -16334
rect 3066 -16570 3072 -16510
rect 3132 -16570 3138 -16510
rect 3072 -16620 3132 -16570
rect 4086 -16620 4146 -16334
rect 4598 -16568 4604 -16508
rect 4664 -16568 4670 -16508
rect 2862 -16626 3132 -16620
rect 3136 -16626 3350 -16620
rect 2862 -16660 2874 -16626
rect 3338 -16660 3350 -16626
rect 2862 -16666 3350 -16660
rect 3880 -16626 4368 -16620
rect 3880 -16660 3892 -16626
rect 4356 -16660 4368 -16626
rect 3880 -16666 4368 -16660
rect 4604 -16710 4664 -16568
rect 5102 -16620 5162 -16142
rect 5620 -16170 5680 -16052
rect 6634 -16052 6654 -15988
rect 6688 -15510 6704 -15476
rect 7656 -15476 7716 -15234
rect 8164 -15386 8224 -15128
rect 7954 -15392 8158 -15386
rect 8164 -15392 8442 -15386
rect 7954 -15426 7966 -15392
rect 8430 -15426 8442 -15392
rect 7954 -15432 8442 -15426
rect 8676 -15476 8736 -15018
rect 9190 -15068 9250 -14910
rect 9696 -15028 9756 -14820
rect 10708 -14820 10726 -14744
rect 10760 -14312 10770 -14244
rect 10760 -14744 10766 -14312
rect 10760 -14820 10768 -14744
rect 11738 -14758 11744 -14320
rect 11732 -14760 11744 -14758
rect 9990 -14870 10478 -14864
rect 9990 -14904 10002 -14870
rect 10466 -14904 10478 -14870
rect 9990 -14910 10478 -14904
rect 9184 -15128 9190 -15068
rect 9250 -15128 9256 -15068
rect 9696 -15088 9922 -15028
rect 10210 -15068 10270 -14910
rect 10708 -14958 10768 -14820
rect 11730 -14820 11744 -14760
rect 12750 -14312 12762 -14244
rect 11778 -14758 11784 -14320
rect 12756 -14754 12762 -14312
rect 11778 -14820 11792 -14758
rect 12744 -14820 12762 -14754
rect 12796 -14312 12810 -14244
rect 13764 -14278 13780 -14244
rect 12796 -14754 12802 -14312
rect 12796 -14820 12804 -14754
rect 13774 -14772 13780 -14278
rect 11008 -14870 11496 -14864
rect 11008 -14904 11020 -14870
rect 11484 -14904 11496 -14870
rect 11008 -14910 11496 -14904
rect 10702 -15018 10708 -14958
rect 10768 -15018 10774 -14958
rect 9190 -15386 9250 -15128
rect 9690 -15234 9696 -15174
rect 9756 -15234 9762 -15174
rect 8972 -15392 9460 -15386
rect 8972 -15426 8984 -15392
rect 9448 -15426 9460 -15392
rect 8972 -15432 9460 -15426
rect 9696 -15476 9756 -15234
rect 9862 -15280 9922 -15088
rect 10204 -15128 10210 -15068
rect 10270 -15128 10276 -15068
rect 9856 -15340 9862 -15280
rect 9922 -15340 9928 -15280
rect 10210 -15386 10270 -15128
rect 9990 -15392 10478 -15386
rect 9990 -15426 10002 -15392
rect 10466 -15426 10478 -15392
rect 9990 -15432 10478 -15426
rect 6688 -15540 6702 -15510
rect 7656 -15520 7672 -15476
rect 6688 -16052 6694 -15540
rect 5918 -16102 6120 -16096
rect 6122 -16102 6406 -16096
rect 5918 -16136 5930 -16102
rect 6394 -16136 6406 -16102
rect 5918 -16142 6120 -16136
rect 6122 -16142 6406 -16136
rect 5614 -16230 5620 -16170
rect 5680 -16230 5686 -16170
rect 5616 -16334 5622 -16274
rect 5682 -16334 5688 -16274
rect 4898 -16626 5386 -16620
rect 4898 -16660 4910 -16626
rect 5374 -16660 5386 -16626
rect 4898 -16666 5386 -16660
rect 2566 -16766 2580 -16710
rect 2574 -17286 2580 -16798
rect 2614 -16766 2626 -16710
rect 3586 -16742 3598 -16710
rect 2614 -17286 2620 -16798
rect 3592 -17242 3598 -16742
rect 2574 -17298 2620 -17286
rect 3586 -17286 3598 -17242
rect 3632 -16742 3646 -16710
rect 4604 -16736 4616 -16710
rect 3632 -17242 3638 -16742
rect 3632 -17286 3646 -17242
rect 2862 -17336 3350 -17330
rect 2862 -17370 2874 -17336
rect 3338 -17370 3350 -17336
rect 2862 -17376 3350 -17370
rect 3586 -17438 3646 -17286
rect 4610 -17286 4616 -16736
rect 4650 -16736 4664 -16710
rect 5622 -16710 5682 -16334
rect 6122 -16620 6182 -16142
rect 6634 -16274 6694 -16052
rect 7666 -16052 7672 -15520
rect 7706 -15510 7718 -15476
rect 7706 -15520 7716 -15510
rect 8676 -15518 8690 -15476
rect 7706 -16052 7712 -15520
rect 8684 -16010 8690 -15518
rect 8676 -16052 8690 -16010
rect 8724 -15518 8736 -15476
rect 8724 -16010 8730 -15518
rect 9692 -15538 9708 -15476
rect 8724 -16052 8736 -16010
rect 9702 -16052 9708 -15538
rect 9742 -15516 9756 -15476
rect 10708 -15476 10768 -15018
rect 11230 -15068 11290 -14910
rect 11224 -15128 11230 -15068
rect 11290 -15128 11296 -15068
rect 11230 -15386 11290 -15128
rect 11730 -15174 11790 -14820
rect 12026 -14870 12514 -14864
rect 12026 -14904 12038 -14870
rect 12502 -14904 12514 -14870
rect 12026 -14910 12372 -14904
rect 12432 -14910 12514 -14904
rect 12232 -15068 12292 -14910
rect 12744 -14958 12804 -14820
rect 13766 -14820 13780 -14772
rect 13814 -14278 13824 -14244
rect 13814 -14772 13820 -14278
rect 14782 -14298 14798 -14244
rect 14792 -14760 14798 -14298
rect 13814 -14820 13826 -14772
rect 13044 -14870 13532 -14864
rect 13044 -14904 13056 -14870
rect 13520 -14904 13532 -14870
rect 13044 -14910 13380 -14904
rect 13440 -14910 13532 -14904
rect 12738 -15018 12744 -14958
rect 12804 -15018 12810 -14958
rect 12226 -15128 12232 -15068
rect 12292 -15128 12298 -15068
rect 11724 -15234 11730 -15174
rect 11790 -15234 11796 -15174
rect 11724 -15340 11730 -15280
rect 11790 -15340 11796 -15280
rect 11008 -15392 11496 -15386
rect 11008 -15426 11020 -15392
rect 11484 -15426 11496 -15392
rect 11008 -15432 11496 -15426
rect 11730 -15476 11790 -15340
rect 12232 -15386 12292 -15128
rect 12026 -15392 12514 -15386
rect 12026 -15426 12038 -15392
rect 12502 -15426 12514 -15392
rect 12026 -15432 12514 -15426
rect 12744 -15476 12804 -15018
rect 13258 -15068 13318 -14910
rect 13252 -15128 13258 -15068
rect 13318 -15128 13324 -15068
rect 13258 -15386 13318 -15128
rect 13766 -15174 13826 -14820
rect 14780 -14820 14798 -14760
rect 14832 -14298 14842 -14244
rect 15802 -14284 15816 -14244
rect 14832 -14760 14838 -14298
rect 15810 -14754 15816 -14284
rect 14832 -14820 14840 -14760
rect 15806 -14780 15816 -14754
rect 14062 -14870 14422 -14864
rect 14482 -14870 14550 -14864
rect 14062 -14904 14074 -14870
rect 14538 -14904 14550 -14870
rect 14062 -14910 14422 -14904
rect 14482 -14910 14550 -14904
rect 14276 -15068 14336 -14910
rect 14780 -14958 14840 -14820
rect 15804 -14820 15816 -14780
rect 15850 -14284 15862 -14244
rect 15850 -14754 15856 -14284
rect 16822 -14298 16834 -14244
rect 15850 -14820 15866 -14754
rect 16828 -14770 16834 -14298
rect 16818 -14820 16834 -14770
rect 16868 -14298 16882 -14244
rect 17844 -14244 17904 -14096
rect 18342 -14160 18402 -13986
rect 16868 -14770 16874 -14298
rect 17844 -14308 17852 -14244
rect 17846 -14764 17852 -14308
rect 16868 -14820 16878 -14770
rect 17838 -14820 17852 -14764
rect 17886 -14308 17904 -14244
rect 18858 -14244 18918 -13854
rect 19362 -13920 19422 -13914
rect 20376 -13920 20436 -13914
rect 19422 -13980 19424 -13974
rect 19362 -13986 19424 -13980
rect 20436 -13980 20438 -13974
rect 20376 -13986 20438 -13980
rect 19364 -14160 19424 -13986
rect 20378 -14160 20438 -13986
rect 20892 -14244 20952 -13854
rect 21400 -13920 21460 -13914
rect 21398 -13980 21400 -13974
rect 21398 -13986 21460 -13980
rect 21398 -14160 21458 -13986
rect 21910 -14096 21916 -14036
rect 21976 -14096 21982 -14036
rect 23042 -14096 23048 -14036
rect 23108 -14096 23114 -14036
rect 21916 -14244 21976 -14096
rect 22206 -14160 22420 -14154
rect 22490 -14160 22694 -14154
rect 22206 -14194 22218 -14160
rect 22682 -14194 22694 -14160
rect 22206 -14200 22694 -14194
rect 18858 -14304 18870 -14244
rect 17886 -14764 17892 -14308
rect 17886 -14766 17898 -14764
rect 17886 -14820 17900 -14766
rect 18864 -14784 18870 -14304
rect 18856 -14820 18870 -14784
rect 18904 -14304 18918 -14244
rect 19874 -14284 19888 -14244
rect 18904 -14784 18910 -14304
rect 19882 -14764 19888 -14284
rect 18904 -14820 18916 -14784
rect 15080 -14870 15568 -14864
rect 15080 -14904 15092 -14870
rect 15556 -14904 15568 -14870
rect 15080 -14910 15568 -14904
rect 14774 -15018 14780 -14958
rect 14840 -15018 14846 -14958
rect 14270 -15128 14276 -15068
rect 14336 -15128 14342 -15068
rect 13760 -15234 13766 -15174
rect 13826 -15234 13832 -15174
rect 13762 -15340 13768 -15280
rect 13828 -15340 13834 -15280
rect 13044 -15392 13532 -15386
rect 13044 -15426 13056 -15392
rect 13520 -15426 13532 -15392
rect 13044 -15432 13532 -15426
rect 13768 -15476 13828 -15340
rect 14276 -15386 14336 -15128
rect 14062 -15392 14550 -15386
rect 14062 -15426 14074 -15392
rect 14538 -15426 14550 -15392
rect 14062 -15432 14550 -15426
rect 14780 -15476 14840 -15018
rect 15284 -15068 15344 -14910
rect 15804 -15036 15864 -14820
rect 16296 -14864 16356 -14862
rect 16098 -14870 16586 -14864
rect 16098 -14904 16110 -14870
rect 16574 -14904 16586 -14870
rect 16098 -14910 16586 -14904
rect 15278 -15128 15284 -15068
rect 15344 -15128 15350 -15068
rect 15648 -15096 15864 -15036
rect 16296 -15068 16356 -14910
rect 16818 -14958 16878 -14820
rect 17328 -14864 17388 -14862
rect 17116 -14870 17604 -14864
rect 17116 -14904 17128 -14870
rect 17592 -14904 17604 -14870
rect 17116 -14910 17604 -14904
rect 18134 -14870 18622 -14864
rect 18134 -14904 18146 -14870
rect 18610 -14904 18622 -14870
rect 18134 -14910 18622 -14904
rect 16812 -15018 16818 -14958
rect 16878 -15018 16884 -14958
rect 15284 -15386 15344 -15128
rect 15648 -15280 15708 -15096
rect 16290 -15128 16296 -15068
rect 16356 -15128 16362 -15068
rect 15796 -15234 15802 -15174
rect 15862 -15234 15868 -15174
rect 15642 -15340 15648 -15280
rect 15708 -15340 15714 -15280
rect 15080 -15392 15568 -15386
rect 15080 -15426 15092 -15392
rect 15556 -15426 15568 -15392
rect 15080 -15432 15568 -15426
rect 9742 -15538 9752 -15516
rect 10708 -15532 10726 -15476
rect 9742 -16052 9748 -15538
rect 10720 -16010 10726 -15532
rect 7666 -16064 7712 -16052
rect 9702 -16064 9748 -16052
rect 10712 -16052 10726 -16010
rect 10760 -15532 10768 -15476
rect 11728 -15528 11744 -15476
rect 10760 -16010 10766 -15532
rect 11738 -15928 11744 -15528
rect 10760 -16052 10772 -16010
rect 11778 -15520 11792 -15476
rect 11778 -15528 11788 -15520
rect 12744 -15524 12762 -15476
rect 11778 -15928 11784 -15528
rect 12756 -16004 12762 -15524
rect 12750 -16052 12762 -16004
rect 12796 -15524 12804 -15476
rect 13764 -15516 13780 -15476
rect 12796 -16004 12802 -15524
rect 13774 -15938 13780 -15516
rect 12796 -16052 12810 -16004
rect 13814 -15514 13830 -15476
rect 13814 -15516 13828 -15514
rect 13814 -15938 13820 -15516
rect 14780 -15522 14798 -15476
rect 14792 -15998 14798 -15522
rect 14780 -16052 14798 -15998
rect 14832 -15522 14840 -15476
rect 15802 -15476 15862 -15234
rect 16296 -15386 16356 -15128
rect 16098 -15392 16586 -15386
rect 16098 -15426 16110 -15392
rect 16574 -15426 16586 -15392
rect 16098 -15432 16586 -15426
rect 16818 -15476 16878 -15018
rect 17328 -15068 17388 -14910
rect 18342 -15068 18402 -14910
rect 18856 -14958 18916 -14820
rect 19872 -14820 19888 -14764
rect 19922 -14284 19934 -14244
rect 19922 -14764 19928 -14284
rect 19922 -14820 19932 -14764
rect 19152 -14870 19640 -14864
rect 19152 -14904 19164 -14870
rect 19628 -14904 19640 -14870
rect 19152 -14910 19420 -14904
rect 19424 -14910 19640 -14904
rect 18850 -15018 18856 -14958
rect 18916 -15018 18922 -14958
rect 17322 -15128 17328 -15068
rect 17388 -15128 17394 -15068
rect 18336 -15128 18342 -15068
rect 18402 -15128 18408 -15068
rect 17328 -15386 17388 -15128
rect 17836 -15234 17842 -15174
rect 17902 -15234 17908 -15174
rect 17116 -15392 17314 -15386
rect 17328 -15392 17604 -15386
rect 17116 -15426 17128 -15392
rect 17592 -15426 17604 -15392
rect 17116 -15432 17604 -15426
rect 17842 -15476 17902 -15234
rect 18342 -15386 18402 -15128
rect 18134 -15392 18402 -15386
rect 18412 -15392 18622 -15386
rect 18134 -15426 18146 -15392
rect 18610 -15426 18622 -15392
rect 18134 -15432 18622 -15426
rect 14832 -15998 14838 -15522
rect 15802 -15528 15816 -15476
rect 14832 -16052 14840 -15998
rect 15810 -16052 15816 -15528
rect 15850 -15518 15866 -15476
rect 15850 -15528 15862 -15518
rect 15850 -16052 15856 -15528
rect 6936 -16102 7424 -16096
rect 6936 -16136 6948 -16102
rect 7412 -16136 7424 -16102
rect 6936 -16142 7132 -16136
rect 7134 -16142 7424 -16136
rect 7954 -16102 8442 -16096
rect 7954 -16136 7966 -16102
rect 8430 -16136 8442 -16102
rect 7954 -16142 8442 -16136
rect 8972 -16102 9460 -16096
rect 8972 -16136 8984 -16102
rect 9448 -16136 9460 -16102
rect 8972 -16142 9460 -16136
rect 9990 -16102 10478 -16096
rect 9990 -16136 10002 -16102
rect 10466 -16136 10478 -16102
rect 9990 -16142 10478 -16136
rect 6628 -16334 6634 -16274
rect 6694 -16334 6700 -16274
rect 6634 -16568 6640 -16508
rect 6700 -16568 6706 -16508
rect 5916 -16626 6120 -16620
rect 6122 -16626 6404 -16620
rect 5916 -16660 5928 -16626
rect 6392 -16660 6404 -16626
rect 5916 -16666 6404 -16660
rect 4650 -17286 4656 -16736
rect 5622 -16742 5634 -16710
rect 5628 -17246 5634 -16742
rect 4610 -17298 4656 -17286
rect 5620 -17286 5634 -17246
rect 5668 -16742 5682 -16710
rect 6640 -16710 6700 -16568
rect 7134 -16620 7194 -16142
rect 7648 -16334 7654 -16274
rect 7714 -16334 7720 -16274
rect 6934 -16626 7132 -16620
rect 7134 -16626 7422 -16620
rect 6934 -16660 6946 -16626
rect 7410 -16660 7422 -16626
rect 6934 -16666 7422 -16660
rect 6640 -16740 6652 -16710
rect 5668 -17246 5674 -16742
rect 5668 -17286 5680 -17246
rect 3880 -17336 4368 -17330
rect 3880 -17370 3892 -17336
rect 4356 -17370 4368 -17336
rect 3880 -17376 4368 -17370
rect 4898 -17336 5386 -17330
rect 4898 -17370 4910 -17336
rect 5374 -17370 5386 -17336
rect 4898 -17376 5386 -17370
rect 2442 -17498 2448 -17438
rect 2508 -17498 2514 -17438
rect 3580 -17498 3586 -17438
rect 3646 -17498 3652 -17438
rect 2330 -17698 2336 -17638
rect 2396 -17698 2402 -17638
rect 2224 -17800 2230 -17740
rect 2290 -17800 2296 -17740
rect 2114 -21252 2120 -21192
rect 2180 -21252 2186 -21192
rect 2230 -21230 2290 -17800
rect 2336 -18874 2396 -17698
rect 2330 -18934 2336 -18874
rect 2396 -18934 2402 -18874
rect 1882 -21402 1888 -21342
rect 1948 -21402 1954 -21342
rect 2120 -24928 2180 -21252
rect 2224 -21290 2230 -21230
rect 2290 -21290 2296 -21230
rect 2230 -23720 2290 -21290
rect 2336 -23594 2396 -18934
rect 2448 -20212 2508 -17498
rect 3578 -17698 3584 -17638
rect 3644 -17698 3650 -17638
rect 3584 -17742 3644 -17698
rect 2568 -17802 3644 -17742
rect 2568 -17804 3132 -17802
rect 2568 -17944 2628 -17804
rect 3072 -17854 3132 -17804
rect 2862 -17860 3350 -17854
rect 2862 -17894 2874 -17860
rect 3338 -17894 3350 -17860
rect 2862 -17900 3350 -17894
rect 2568 -17976 2580 -17944
rect 2574 -18520 2580 -17976
rect 2614 -17976 2628 -17944
rect 3584 -17944 3644 -17802
rect 4088 -17854 4148 -17376
rect 4596 -17578 4602 -17518
rect 4662 -17578 4668 -17518
rect 3880 -17860 4368 -17854
rect 3880 -17894 3892 -17860
rect 4356 -17894 4368 -17860
rect 3880 -17900 4368 -17894
rect 2614 -18520 2620 -17976
rect 3584 -17980 3598 -17944
rect 2574 -18532 2620 -18520
rect 3592 -18520 3598 -17980
rect 3632 -17980 3644 -17944
rect 4602 -17944 4662 -17578
rect 5116 -17632 5176 -17376
rect 5620 -17414 5680 -17286
rect 6646 -17286 6652 -16740
rect 6686 -16740 6700 -16710
rect 7654 -16710 7714 -16334
rect 8160 -16620 8220 -16142
rect 8670 -16230 8676 -16170
rect 8736 -16230 8742 -16170
rect 7952 -16626 8440 -16620
rect 7952 -16660 7964 -16626
rect 8428 -16660 8440 -16626
rect 7952 -16666 8440 -16660
rect 6686 -17286 6692 -16740
rect 7654 -16754 7670 -16710
rect 7664 -17236 7670 -16754
rect 6646 -17298 6692 -17286
rect 7656 -17286 7670 -17236
rect 7704 -16754 7714 -16710
rect 8676 -16710 8736 -16230
rect 10712 -16274 10772 -16052
rect 11008 -16102 11176 -16096
rect 12424 -16102 12514 -16096
rect 11008 -16136 11020 -16102
rect 12502 -16136 12514 -16102
rect 11008 -16142 11176 -16136
rect 12424 -16142 12514 -16136
rect 12750 -16274 12810 -16052
rect 15810 -16064 15856 -16052
rect 16818 -16052 16834 -15476
rect 16868 -16052 16878 -15476
rect 17838 -15518 17852 -15476
rect 17842 -15538 17852 -15518
rect 13044 -16102 13236 -16096
rect 14480 -16102 14550 -16096
rect 13044 -16136 13056 -16102
rect 14538 -16136 14550 -16102
rect 13044 -16142 13236 -16136
rect 14480 -16142 14550 -16136
rect 15080 -16102 15568 -16096
rect 15080 -16136 15092 -16102
rect 15556 -16136 15568 -16102
rect 15080 -16142 15568 -16136
rect 16098 -16102 16586 -16096
rect 16098 -16136 16110 -16102
rect 16574 -16136 16586 -16102
rect 16098 -16142 16586 -16136
rect 14776 -16230 14782 -16170
rect 14842 -16230 14848 -16170
rect 10706 -16334 10712 -16274
rect 10772 -16334 10778 -16274
rect 12744 -16334 12750 -16274
rect 12810 -16334 12816 -16274
rect 9690 -16456 9696 -16396
rect 9756 -16456 9762 -16396
rect 11724 -16456 11730 -16396
rect 11790 -16456 11796 -16396
rect 13754 -16456 13760 -16396
rect 13820 -16456 13826 -16396
rect 8970 -16626 9458 -16620
rect 8970 -16660 8982 -16626
rect 9446 -16660 9458 -16626
rect 8970 -16666 9458 -16660
rect 7704 -17236 7710 -16754
rect 8676 -16772 8688 -16710
rect 7704 -17286 7716 -17236
rect 8682 -17250 8688 -16772
rect 5916 -17336 6404 -17330
rect 5916 -17370 5928 -17336
rect 6392 -17370 6404 -17336
rect 5916 -17376 6404 -17370
rect 6934 -17336 7422 -17330
rect 6934 -17370 6946 -17336
rect 7410 -17370 7422 -17336
rect 6934 -17376 7422 -17370
rect 5614 -17474 5620 -17414
rect 5680 -17474 5686 -17414
rect 5110 -17692 5116 -17632
rect 5176 -17692 5182 -17632
rect 5116 -17854 5176 -17692
rect 4898 -17860 5386 -17854
rect 4898 -17894 4910 -17860
rect 5374 -17894 5386 -17860
rect 4898 -17900 5386 -17894
rect 3632 -18520 3638 -17980
rect 4602 -17986 4616 -17944
rect 4610 -18462 4616 -17986
rect 3592 -18532 3638 -18520
rect 4604 -18520 4616 -18462
rect 4650 -17986 4662 -17944
rect 5620 -17944 5680 -17474
rect 6118 -17626 6178 -17376
rect 6636 -17578 6642 -17518
rect 6702 -17578 6708 -17518
rect 6118 -17632 6180 -17626
rect 6118 -17692 6120 -17632
rect 6118 -17698 6180 -17692
rect 6118 -17854 6178 -17698
rect 5916 -17860 6404 -17854
rect 5916 -17894 5928 -17860
rect 6392 -17894 6404 -17860
rect 5916 -17900 6404 -17894
rect 4650 -18462 4656 -17986
rect 5620 -17988 5634 -17944
rect 4650 -18520 4664 -18462
rect 5628 -18472 5634 -17988
rect 2862 -18570 3350 -18564
rect 2862 -18604 2874 -18570
rect 3338 -18604 3350 -18570
rect 2862 -18610 3350 -18604
rect 3880 -18570 4368 -18564
rect 3880 -18604 3892 -18570
rect 4356 -18604 4368 -18570
rect 3880 -18610 4368 -18604
rect 3578 -18730 3584 -18670
rect 3644 -18730 3650 -18670
rect 2862 -19092 3350 -19086
rect 2862 -19126 2874 -19092
rect 3338 -19126 3350 -19092
rect 2862 -19132 3350 -19126
rect 2574 -19176 2620 -19164
rect 2574 -19706 2580 -19176
rect 2564 -19752 2580 -19706
rect 2614 -19706 2620 -19176
rect 3584 -19176 3644 -18730
rect 4090 -18772 4150 -18610
rect 4084 -18832 4090 -18772
rect 4150 -18832 4156 -18772
rect 4604 -18974 4664 -18520
rect 5622 -18520 5634 -18472
rect 5668 -17988 5680 -17944
rect 6642 -17944 6702 -17578
rect 7134 -17626 7194 -17376
rect 7656 -17414 7716 -17286
rect 8674 -17286 8688 -17250
rect 8722 -16772 8736 -16710
rect 9696 -16710 9756 -16456
rect 9988 -16626 10476 -16620
rect 9988 -16660 10000 -16626
rect 10464 -16660 10476 -16626
rect 9988 -16666 10476 -16660
rect 11006 -16626 11494 -16620
rect 11006 -16660 11018 -16626
rect 11482 -16660 11494 -16626
rect 11006 -16666 11494 -16660
rect 9696 -16766 9706 -16710
rect 8722 -17250 8728 -16772
rect 8722 -17286 8734 -17250
rect 7952 -17336 8440 -17330
rect 7952 -17370 7964 -17336
rect 8428 -17370 8440 -17336
rect 7952 -17376 8440 -17370
rect 7650 -17474 7656 -17414
rect 7716 -17474 7722 -17414
rect 7132 -17632 7194 -17626
rect 7192 -17692 7194 -17632
rect 7132 -17698 7194 -17692
rect 7134 -17854 7194 -17698
rect 6934 -17860 7422 -17854
rect 6934 -17894 6946 -17860
rect 7410 -17894 7422 -17860
rect 6934 -17900 7422 -17894
rect 6642 -17986 6652 -17944
rect 5668 -18472 5674 -17988
rect 5668 -18520 5682 -18472
rect 4898 -18570 5386 -18564
rect 4898 -18604 4910 -18570
rect 5374 -18604 5386 -18570
rect 4898 -18610 5386 -18604
rect 5622 -18670 5682 -18520
rect 6646 -18520 6652 -17986
rect 6686 -17986 6702 -17944
rect 7656 -17944 7716 -17474
rect 8152 -17632 8212 -17376
rect 8674 -17518 8734 -17286
rect 9700 -17286 9706 -16766
rect 9740 -16766 9756 -16710
rect 10718 -16710 10764 -16698
rect 9740 -17286 9746 -16766
rect 10718 -17256 10724 -16710
rect 9700 -17298 9746 -17286
rect 10708 -17286 10724 -17256
rect 10758 -17256 10764 -16710
rect 11730 -16710 11790 -16456
rect 12024 -16626 12512 -16620
rect 12024 -16660 12036 -16626
rect 12500 -16660 12512 -16626
rect 12024 -16666 12512 -16660
rect 13042 -16626 13530 -16620
rect 13042 -16660 13054 -16626
rect 13518 -16660 13530 -16626
rect 13042 -16666 13530 -16660
rect 11730 -16760 11742 -16710
rect 10758 -17286 10768 -17256
rect 8970 -17336 9458 -17330
rect 8970 -17370 8982 -17336
rect 9446 -17370 9458 -17336
rect 8970 -17376 9458 -17370
rect 9988 -17336 10476 -17330
rect 9988 -17370 10000 -17336
rect 10464 -17370 10476 -17336
rect 9988 -17376 10476 -17370
rect 8668 -17578 8674 -17518
rect 8734 -17578 8740 -17518
rect 9164 -17574 9224 -17376
rect 10206 -17574 10266 -17376
rect 10708 -17518 10768 -17286
rect 11736 -17286 11742 -16760
rect 11776 -16760 11790 -16710
rect 12754 -16710 12800 -16698
rect 11776 -17286 11782 -16760
rect 12754 -17244 12760 -16710
rect 11736 -17298 11782 -17286
rect 12748 -17286 12760 -17244
rect 12794 -17244 12800 -16710
rect 13760 -16710 13820 -16456
rect 14060 -16626 14548 -16620
rect 14060 -16660 14072 -16626
rect 14536 -16660 14548 -16626
rect 14060 -16666 14548 -16660
rect 13760 -16754 13778 -16710
rect 12794 -17286 12808 -17244
rect 11006 -17336 11494 -17330
rect 11006 -17370 11018 -17336
rect 11482 -17370 11494 -17336
rect 11006 -17376 11494 -17370
rect 12024 -17336 12512 -17330
rect 12024 -17370 12036 -17336
rect 12500 -17370 12512 -17336
rect 12024 -17376 12512 -17370
rect 8668 -17690 8674 -17630
rect 8734 -17690 8740 -17630
rect 9164 -17634 10266 -17574
rect 10702 -17578 10708 -17518
rect 10768 -17578 10774 -17518
rect 8152 -17854 8212 -17692
rect 7952 -17860 8440 -17854
rect 7952 -17894 7964 -17860
rect 8428 -17894 8440 -17860
rect 7952 -17900 8440 -17894
rect 6686 -18520 6692 -17986
rect 7656 -17992 7670 -17944
rect 7664 -18470 7670 -17992
rect 6646 -18532 6692 -18520
rect 7658 -18520 7670 -18470
rect 7704 -17992 7716 -17944
rect 8674 -17944 8734 -17690
rect 9164 -17854 9224 -17634
rect 9686 -17800 9692 -17740
rect 9752 -17800 9758 -17740
rect 8970 -17860 9458 -17854
rect 8970 -17894 8982 -17860
rect 9446 -17894 9458 -17860
rect 8970 -17900 9458 -17894
rect 7704 -18470 7710 -17992
rect 8674 -18002 8688 -17944
rect 7704 -18520 7718 -18470
rect 5916 -18570 6404 -18564
rect 5916 -18604 5928 -18570
rect 6392 -18604 6404 -18570
rect 5916 -18610 6404 -18604
rect 6934 -18570 7422 -18564
rect 6934 -18604 6946 -18570
rect 7410 -18604 7422 -18570
rect 6934 -18610 7422 -18604
rect 5616 -18730 5622 -18670
rect 5682 -18730 5688 -18670
rect 5614 -18934 5620 -18874
rect 5680 -18934 5686 -18874
rect 6128 -18880 6188 -18610
rect 7150 -18880 7210 -18610
rect 7658 -18670 7718 -18520
rect 8682 -18520 8688 -18002
rect 8722 -18002 8734 -17944
rect 9692 -17944 9752 -17800
rect 10206 -17854 10266 -17634
rect 10704 -17690 10710 -17630
rect 10770 -17690 10776 -17630
rect 9988 -17860 10476 -17854
rect 9988 -17894 10000 -17860
rect 10464 -17894 10476 -17860
rect 9988 -17900 10476 -17894
rect 9692 -17990 9706 -17944
rect 8722 -18520 8728 -18002
rect 8682 -18532 8728 -18520
rect 9700 -18520 9706 -17990
rect 9740 -17990 9752 -17944
rect 10710 -17944 10770 -17690
rect 11206 -17854 11266 -17376
rect 11720 -17800 11726 -17740
rect 11786 -17800 11792 -17740
rect 11006 -17860 11494 -17854
rect 11006 -17894 11018 -17860
rect 11482 -17894 11494 -17860
rect 11006 -17900 11494 -17894
rect 9740 -18520 9746 -17990
rect 10710 -18012 10724 -17944
rect 9700 -18532 9746 -18520
rect 10718 -18520 10724 -18012
rect 10758 -18012 10770 -17944
rect 11726 -17944 11786 -17800
rect 12240 -17854 12300 -17376
rect 12748 -17518 12808 -17286
rect 13772 -17286 13778 -16754
rect 13812 -16754 13820 -16710
rect 14782 -16710 14842 -16230
rect 15304 -16620 15364 -16142
rect 15794 -16334 15800 -16274
rect 15860 -16334 15866 -16274
rect 15078 -16626 15566 -16620
rect 15078 -16660 15090 -16626
rect 15554 -16660 15566 -16626
rect 15078 -16666 15566 -16660
rect 13812 -17286 13818 -16754
rect 14782 -16762 14796 -16710
rect 14790 -17234 14796 -16762
rect 13772 -17298 13818 -17286
rect 14782 -17286 14796 -17234
rect 14830 -16762 14842 -16710
rect 15800 -16710 15860 -16334
rect 16306 -16620 16366 -16142
rect 16818 -16274 16878 -16052
rect 17846 -16052 17852 -15538
rect 17886 -15538 17902 -15476
rect 18856 -15476 18916 -15018
rect 19360 -15068 19420 -14910
rect 19354 -15128 19360 -15068
rect 19420 -15128 19426 -15068
rect 19360 -15386 19420 -15128
rect 19872 -15174 19932 -14820
rect 20892 -14820 20906 -14244
rect 20940 -14276 20954 -14244
rect 21912 -14272 21924 -14244
rect 20940 -14820 20952 -14276
rect 21916 -14308 21924 -14272
rect 21918 -14760 21924 -14308
rect 20170 -14870 20658 -14864
rect 20170 -14904 20182 -14870
rect 20646 -14904 20658 -14870
rect 20170 -14910 20658 -14904
rect 20384 -15068 20444 -14910
rect 20892 -14958 20952 -14820
rect 21912 -14820 21924 -14760
rect 21958 -14308 21976 -14244
rect 21958 -14760 21964 -14308
rect 21958 -14820 21972 -14760
rect 22936 -14772 22942 -14284
rect 21188 -14870 21676 -14864
rect 21188 -14904 21200 -14870
rect 21664 -14904 21676 -14870
rect 21188 -14910 21676 -14904
rect 20886 -15018 20892 -14958
rect 20952 -15018 20958 -14958
rect 20378 -15128 20384 -15068
rect 20444 -15128 20450 -15068
rect 19866 -15234 19872 -15174
rect 19932 -15234 19938 -15174
rect 19866 -15338 19872 -15278
rect 19932 -15338 19938 -15278
rect 19152 -15392 19352 -15386
rect 19360 -15392 19640 -15386
rect 19152 -15426 19164 -15392
rect 19628 -15426 19640 -15392
rect 19152 -15432 19640 -15426
rect 19352 -15444 19412 -15432
rect 19872 -15476 19932 -15338
rect 20384 -15386 20444 -15128
rect 20170 -15392 20658 -15386
rect 20170 -15426 20182 -15392
rect 20646 -15426 20658 -15392
rect 20170 -15432 20658 -15426
rect 18856 -15534 18870 -15476
rect 17886 -16052 17892 -15538
rect 18864 -16004 18870 -15534
rect 17846 -16064 17892 -16052
rect 18854 -16052 18870 -16004
rect 18904 -15534 18916 -15476
rect 19870 -15522 19888 -15476
rect 18904 -16004 18910 -15534
rect 19872 -15550 19888 -15522
rect 19882 -15998 19888 -15550
rect 18904 -16052 18914 -16004
rect 17116 -16102 17604 -16096
rect 17116 -16136 17128 -16102
rect 17318 -16136 17378 -16134
rect 17592 -16136 17604 -16102
rect 17116 -16142 17604 -16136
rect 18134 -16102 18622 -16096
rect 18134 -16136 18146 -16102
rect 18352 -16136 18412 -16130
rect 18610 -16136 18622 -16102
rect 18134 -16142 18622 -16136
rect 16812 -16334 16818 -16274
rect 16878 -16334 16884 -16274
rect 17318 -16620 17378 -16142
rect 17832 -16334 17838 -16274
rect 17898 -16334 17904 -16274
rect 16096 -16626 16584 -16620
rect 16096 -16660 16108 -16626
rect 16572 -16660 16584 -16626
rect 16096 -16666 16584 -16660
rect 17114 -16626 17602 -16620
rect 17114 -16660 17126 -16626
rect 17590 -16660 17602 -16626
rect 17114 -16666 17602 -16660
rect 15800 -16758 15814 -16710
rect 14830 -17234 14836 -16762
rect 14830 -17286 14842 -17234
rect 15808 -17254 15814 -16758
rect 13042 -17336 13530 -17330
rect 13042 -17370 13054 -17336
rect 13518 -17370 13530 -17336
rect 13042 -17376 13530 -17370
rect 14060 -17336 14548 -17330
rect 14060 -17370 14072 -17336
rect 14536 -17370 14548 -17336
rect 14060 -17376 14548 -17370
rect 12742 -17578 12748 -17518
rect 12808 -17578 12814 -17518
rect 13262 -17574 13322 -17376
rect 14270 -17574 14330 -17376
rect 14782 -17518 14842 -17286
rect 15800 -17286 15814 -17254
rect 15848 -16758 15860 -16710
rect 16826 -16710 16872 -16698
rect 15848 -17254 15854 -16758
rect 16826 -17250 16832 -16710
rect 15848 -17286 15860 -17254
rect 15078 -17336 15566 -17330
rect 15078 -17370 15090 -17336
rect 15554 -17370 15566 -17336
rect 15078 -17376 15566 -17370
rect 12740 -17690 12746 -17630
rect 12806 -17690 12812 -17630
rect 13262 -17634 14330 -17574
rect 14776 -17578 14782 -17518
rect 14842 -17578 14848 -17518
rect 14972 -17582 14978 -17522
rect 15038 -17582 15044 -17522
rect 12024 -17860 12512 -17854
rect 12024 -17894 12036 -17860
rect 12500 -17894 12512 -17860
rect 12024 -17900 12512 -17894
rect 11726 -17992 11742 -17944
rect 10758 -18520 10764 -18012
rect 10718 -18532 10764 -18520
rect 11736 -18520 11742 -17992
rect 11776 -17992 11786 -17944
rect 12746 -17944 12806 -17690
rect 13262 -17854 13322 -17634
rect 13760 -17800 13766 -17740
rect 13826 -17800 13832 -17740
rect 13042 -17860 13530 -17854
rect 13042 -17894 13054 -17860
rect 13518 -17894 13530 -17860
rect 13042 -17900 13530 -17894
rect 11776 -18520 11782 -17992
rect 12746 -17994 12760 -17944
rect 11736 -18532 11782 -18520
rect 12754 -18520 12760 -17994
rect 12794 -17994 12806 -17944
rect 13766 -17944 13826 -17800
rect 14270 -17854 14330 -17634
rect 14776 -17690 14782 -17630
rect 14842 -17690 14848 -17630
rect 14060 -17860 14548 -17854
rect 14060 -17894 14072 -17860
rect 14536 -17894 14548 -17860
rect 14060 -17900 14548 -17894
rect 13766 -17982 13778 -17944
rect 12794 -18520 12800 -17994
rect 13772 -18474 13778 -17982
rect 12754 -18532 12800 -18520
rect 13766 -18520 13778 -18474
rect 13812 -17982 13826 -17944
rect 14782 -17944 14842 -17690
rect 14978 -17740 15038 -17582
rect 15272 -17738 15332 -17376
rect 15800 -17414 15860 -17286
rect 16816 -17286 16832 -17250
rect 16866 -17250 16872 -16710
rect 17838 -16710 17898 -16334
rect 18352 -16620 18412 -16142
rect 18854 -16274 18914 -16052
rect 19876 -16052 19888 -15998
rect 19922 -15550 19932 -15476
rect 20892 -15476 20952 -15018
rect 21404 -15068 21464 -14910
rect 21912 -14968 21972 -14820
rect 22928 -14820 22942 -14772
rect 22976 -14772 22982 -14284
rect 22976 -14820 22988 -14772
rect 22206 -14870 22694 -14864
rect 22206 -14904 22218 -14870
rect 22682 -14904 22694 -14870
rect 22206 -14910 22694 -14904
rect 22422 -14968 22482 -14910
rect 22928 -14968 22988 -14820
rect 23048 -14968 23108 -14096
rect 21912 -15028 23108 -14968
rect 21398 -15128 21404 -15068
rect 21464 -15128 21470 -15068
rect 21404 -15386 21464 -15128
rect 21906 -15234 21912 -15174
rect 21972 -15234 21978 -15174
rect 21912 -15276 21972 -15234
rect 21912 -15336 22990 -15276
rect 23048 -15278 23108 -15028
rect 21188 -15392 21676 -15386
rect 21188 -15426 21200 -15392
rect 21664 -15426 21676 -15392
rect 21188 -15432 21676 -15426
rect 20892 -15502 20906 -15476
rect 19922 -15998 19928 -15550
rect 20900 -15994 20906 -15502
rect 19922 -16052 19936 -15998
rect 19152 -16102 19640 -16096
rect 19152 -16136 19164 -16102
rect 19628 -16136 19640 -16102
rect 19152 -16142 19368 -16136
rect 19428 -16142 19640 -16136
rect 19876 -16170 19936 -16052
rect 20890 -16052 20906 -15994
rect 20940 -15502 20952 -15476
rect 21912 -15476 21972 -15336
rect 22398 -15386 22458 -15336
rect 22206 -15392 22458 -15386
rect 22476 -15392 22694 -15386
rect 22206 -15426 22218 -15392
rect 22682 -15426 22694 -15392
rect 22206 -15432 22694 -15426
rect 22930 -15476 22990 -15336
rect 23042 -15338 23048 -15278
rect 23108 -15338 23114 -15278
rect 20940 -15994 20946 -15502
rect 21912 -15532 21924 -15476
rect 20940 -16052 20950 -15994
rect 20170 -16102 20658 -16096
rect 20170 -16136 20182 -16102
rect 20646 -16136 20658 -16102
rect 20170 -16142 20658 -16136
rect 19870 -16230 19876 -16170
rect 19936 -16230 19942 -16170
rect 20890 -16274 20950 -16052
rect 21918 -16052 21924 -15532
rect 21958 -15532 21972 -15476
rect 22926 -15512 22942 -15476
rect 22930 -15518 22942 -15512
rect 21958 -16052 21964 -15532
rect 22936 -15970 22942 -15518
rect 21918 -16064 21964 -16052
rect 22932 -16052 22942 -16008
rect 22976 -15518 22990 -15476
rect 22976 -15970 22982 -15518
rect 22976 -16052 22992 -16008
rect 21188 -16102 21676 -16096
rect 21188 -16136 21200 -16102
rect 21664 -16136 21676 -16102
rect 21188 -16142 21676 -16136
rect 22206 -16102 22694 -16096
rect 22206 -16136 22218 -16102
rect 22682 -16136 22694 -16102
rect 22206 -16142 22694 -16136
rect 18848 -16334 18854 -16274
rect 18914 -16334 18920 -16274
rect 20884 -16334 20890 -16274
rect 20950 -16334 20956 -16274
rect 21380 -16620 21440 -16142
rect 22932 -16178 22992 -16052
rect 22932 -16238 23222 -16178
rect 22418 -16544 22986 -16484
rect 22418 -16620 22478 -16544
rect 18132 -16626 18620 -16620
rect 18132 -16660 18144 -16626
rect 18608 -16660 18620 -16626
rect 18132 -16666 18620 -16660
rect 19150 -16626 19638 -16620
rect 19150 -16660 19162 -16626
rect 19626 -16660 19638 -16626
rect 19150 -16666 19638 -16660
rect 20168 -16626 20656 -16620
rect 20168 -16660 20180 -16626
rect 20644 -16660 20656 -16626
rect 20168 -16666 20656 -16660
rect 21186 -16626 21674 -16620
rect 21186 -16660 21198 -16626
rect 21662 -16660 21674 -16626
rect 21186 -16666 21674 -16660
rect 22204 -16626 22692 -16620
rect 22204 -16660 22216 -16626
rect 22680 -16660 22692 -16626
rect 22204 -16666 22692 -16660
rect 17838 -16768 17850 -16710
rect 17844 -17240 17850 -16768
rect 16866 -17286 16876 -17250
rect 16096 -17336 16584 -17330
rect 16096 -17370 16108 -17336
rect 16572 -17370 16584 -17336
rect 16096 -17376 16584 -17370
rect 15794 -17474 15800 -17414
rect 15860 -17474 15866 -17414
rect 14972 -17800 14978 -17740
rect 15038 -17800 15044 -17740
rect 15266 -17798 15272 -17738
rect 15332 -17798 15338 -17738
rect 15272 -17854 15332 -17798
rect 15078 -17860 15566 -17854
rect 15078 -17894 15090 -17860
rect 15554 -17894 15566 -17860
rect 15078 -17900 15566 -17894
rect 13812 -18474 13818 -17982
rect 14782 -17988 14796 -17944
rect 13812 -18520 13826 -18474
rect 7952 -18570 8440 -18564
rect 7952 -18604 7964 -18570
rect 8428 -18604 8440 -18570
rect 7952 -18610 8440 -18604
rect 8970 -18570 9458 -18564
rect 8970 -18604 8982 -18570
rect 9446 -18604 9458 -18570
rect 8970 -18610 9458 -18604
rect 9988 -18570 10476 -18564
rect 9988 -18604 10000 -18570
rect 10464 -18604 10476 -18570
rect 9988 -18610 10476 -18604
rect 11006 -18570 11494 -18564
rect 11006 -18604 11018 -18570
rect 11482 -18604 11494 -18570
rect 11006 -18610 11494 -18604
rect 12024 -18570 12512 -18564
rect 12024 -18604 12036 -18570
rect 12500 -18604 12512 -18570
rect 12024 -18610 12238 -18604
rect 12240 -18610 12512 -18604
rect 13042 -18570 13530 -18564
rect 13042 -18604 13054 -18570
rect 13518 -18604 13530 -18570
rect 13042 -18610 13264 -18604
rect 13268 -18610 13530 -18604
rect 7652 -18730 7658 -18670
rect 7718 -18730 7724 -18670
rect 4598 -19034 4604 -18974
rect 4664 -19034 4670 -18974
rect 3880 -19092 4368 -19086
rect 3880 -19126 3892 -19092
rect 4356 -19126 4368 -19092
rect 3880 -19132 4368 -19126
rect 3584 -19214 3598 -19176
rect 2614 -19752 2624 -19706
rect 3592 -19710 3598 -19214
rect 2564 -19914 2624 -19752
rect 3582 -19752 3598 -19710
rect 3632 -19214 3644 -19176
rect 4604 -19176 4664 -19034
rect 4898 -19092 5386 -19086
rect 4898 -19126 4910 -19092
rect 5374 -19126 5386 -19092
rect 4898 -19132 5386 -19126
rect 3632 -19710 3638 -19214
rect 4604 -19216 4616 -19176
rect 3632 -19752 3642 -19710
rect 2862 -19802 3350 -19796
rect 2862 -19836 2874 -19802
rect 3338 -19836 3350 -19802
rect 2862 -19842 3350 -19836
rect 3076 -19914 3136 -19842
rect 3582 -19914 3642 -19752
rect 4610 -19752 4616 -19216
rect 4650 -19216 4664 -19176
rect 5620 -19176 5680 -18934
rect 6122 -18940 6128 -18880
rect 6188 -18940 6194 -18880
rect 7144 -18940 7150 -18880
rect 7210 -18940 7216 -18880
rect 6632 -19034 6638 -18974
rect 6698 -19034 6704 -18974
rect 5916 -19092 6404 -19086
rect 5916 -19126 5928 -19092
rect 6392 -19126 6404 -19092
rect 5916 -19132 6404 -19126
rect 4650 -19752 4656 -19216
rect 5620 -19228 5634 -19176
rect 4610 -19764 4656 -19752
rect 5628 -19752 5634 -19228
rect 5668 -19228 5680 -19176
rect 6638 -19176 6698 -19034
rect 7150 -19086 7210 -18940
rect 6934 -19092 7422 -19086
rect 6934 -19126 6946 -19092
rect 7410 -19126 7422 -19092
rect 6934 -19132 7422 -19126
rect 6638 -19220 6652 -19176
rect 5668 -19752 5674 -19228
rect 6646 -19716 6652 -19220
rect 5628 -19764 5674 -19752
rect 6638 -19752 6652 -19716
rect 6686 -19220 6698 -19176
rect 7658 -19176 7718 -18730
rect 8164 -18880 8224 -18610
rect 9182 -18772 9242 -18610
rect 10202 -18660 10262 -18610
rect 11202 -18660 11262 -18610
rect 12240 -18660 12300 -18610
rect 13268 -18660 13328 -18610
rect 9684 -18730 9690 -18670
rect 9750 -18730 9756 -18670
rect 10202 -18720 13328 -18660
rect 9176 -18832 9182 -18772
rect 9242 -18832 9248 -18772
rect 8158 -18940 8164 -18880
rect 8224 -18940 8230 -18880
rect 9176 -18940 9182 -18880
rect 9242 -18940 9248 -18880
rect 8164 -19086 8224 -18940
rect 8668 -19034 8674 -18974
rect 8734 -19034 8740 -18974
rect 7952 -19092 8440 -19086
rect 7952 -19126 7964 -19092
rect 8428 -19126 8440 -19092
rect 7952 -19132 8440 -19126
rect 6686 -19716 6692 -19220
rect 6686 -19752 6698 -19716
rect 3880 -19802 4368 -19796
rect 3880 -19836 3892 -19802
rect 4356 -19836 4368 -19802
rect 3880 -19842 4368 -19836
rect 4898 -19802 5386 -19796
rect 4898 -19836 4910 -19802
rect 5374 -19836 5386 -19802
rect 4898 -19842 5386 -19836
rect 5916 -19802 6404 -19796
rect 5916 -19836 5928 -19802
rect 6392 -19836 6404 -19802
rect 5916 -19842 6404 -19836
rect 4086 -19898 4146 -19842
rect 2564 -19974 3642 -19914
rect 4080 -19958 4086 -19898
rect 4146 -19958 4152 -19898
rect 4990 -19958 4996 -19898
rect 5056 -19958 5062 -19898
rect 4080 -20174 4086 -20114
rect 4146 -20174 4152 -20114
rect 4086 -20180 4148 -20174
rect 2448 -20218 2510 -20212
rect 2448 -20278 2450 -20218
rect 2448 -20284 2510 -20278
rect 2448 -22462 2508 -20284
rect 4088 -20320 4148 -20180
rect 4996 -20320 5056 -19958
rect 5124 -20114 5184 -19842
rect 5992 -19958 5998 -19898
rect 6058 -19958 6064 -19898
rect 5124 -20180 5184 -20174
rect 5998 -20320 6058 -19958
rect 6138 -20114 6198 -19842
rect 6638 -20000 6698 -19752
rect 7658 -19752 7670 -19176
rect 7704 -19752 7718 -19176
rect 8674 -19176 8734 -19034
rect 9182 -19086 9242 -18940
rect 8970 -19092 9458 -19086
rect 8970 -19126 8982 -19092
rect 9446 -19126 9458 -19092
rect 8970 -19132 9458 -19126
rect 8674 -19212 8688 -19176
rect 6934 -19802 7422 -19796
rect 6934 -19836 6946 -19802
rect 7410 -19836 7422 -19802
rect 6934 -19842 7126 -19836
rect 7150 -19842 7422 -19836
rect 7150 -19898 7210 -19842
rect 7144 -19958 7150 -19898
rect 7210 -19958 7216 -19898
rect 6632 -20060 6638 -20000
rect 6698 -20060 6704 -20000
rect 6132 -20174 6138 -20114
rect 6198 -20174 6204 -20114
rect 7150 -20320 7210 -19958
rect 2862 -20326 3350 -20320
rect 2862 -20360 2874 -20326
rect 3338 -20360 3350 -20326
rect 2862 -20366 3350 -20360
rect 3880 -20326 4368 -20320
rect 3880 -20360 3892 -20326
rect 4356 -20360 4368 -20326
rect 3880 -20366 4368 -20360
rect 4898 -20326 5386 -20320
rect 4898 -20360 4910 -20326
rect 5374 -20360 5386 -20326
rect 4898 -20366 5386 -20360
rect 5916 -20326 6404 -20320
rect 5916 -20360 5928 -20326
rect 6392 -20360 6404 -20326
rect 5916 -20366 6404 -20360
rect 6934 -20326 7422 -20320
rect 6934 -20360 6946 -20326
rect 7410 -20360 7422 -20326
rect 6934 -20366 7422 -20360
rect 2574 -20410 2620 -20398
rect 2574 -20948 2580 -20410
rect 2568 -20986 2580 -20948
rect 2614 -20948 2620 -20410
rect 3592 -20410 3638 -20398
rect 3592 -20948 3598 -20410
rect 2614 -20986 2628 -20948
rect 2568 -21116 2628 -20986
rect 3586 -20986 3598 -20948
rect 3632 -20948 3638 -20410
rect 4610 -20410 4656 -20398
rect 4610 -20936 4616 -20410
rect 3632 -20986 3646 -20948
rect 2862 -21036 3350 -21030
rect 2862 -21070 2874 -21036
rect 3338 -21070 3350 -21036
rect 2862 -21076 3350 -21070
rect 3066 -21116 3126 -21076
rect 3586 -21116 3646 -20986
rect 4602 -20986 4616 -20936
rect 4650 -20936 4656 -20410
rect 5628 -20410 5674 -20398
rect 5628 -20928 5634 -20410
rect 4650 -20986 4662 -20936
rect 3880 -21036 4368 -21030
rect 3880 -21070 3892 -21036
rect 4356 -21070 4368 -21036
rect 3880 -21076 4368 -21070
rect 2568 -21176 3646 -21116
rect 3586 -21230 3646 -21176
rect 4078 -21186 4084 -21126
rect 4144 -21186 4150 -21126
rect 3580 -21290 3586 -21230
rect 3646 -21290 3652 -21230
rect 3576 -21500 3582 -21440
rect 3642 -21500 3648 -21440
rect 2862 -21560 3350 -21554
rect 2862 -21594 2874 -21560
rect 3338 -21594 3350 -21560
rect 2862 -21600 3350 -21594
rect 2574 -21644 2620 -21632
rect 2574 -22186 2580 -21644
rect 2564 -22220 2580 -22186
rect 2614 -22186 2620 -21644
rect 3582 -21644 3642 -21500
rect 4084 -21554 4144 -21186
rect 4602 -21342 4662 -20986
rect 5620 -20986 5634 -20928
rect 5668 -20928 5674 -20410
rect 6646 -20410 6692 -20398
rect 5668 -20986 5680 -20928
rect 6646 -20940 6652 -20410
rect 4898 -21036 5386 -21030
rect 4898 -21070 4910 -21036
rect 5374 -21070 5386 -21036
rect 4898 -21076 5386 -21070
rect 5092 -21126 5152 -21076
rect 5086 -21186 5092 -21126
rect 5152 -21186 5158 -21126
rect 4596 -21402 4602 -21342
rect 4662 -21402 4668 -21342
rect 5620 -21440 5680 -20986
rect 6640 -20986 6652 -20940
rect 6686 -20940 6692 -20410
rect 7658 -20410 7718 -19752
rect 8682 -19752 8688 -19212
rect 8722 -19212 8734 -19176
rect 9690 -19176 9750 -18730
rect 10196 -18940 10202 -18880
rect 10262 -18940 10268 -18880
rect 13268 -18896 13328 -18720
rect 13766 -18786 13826 -18520
rect 14790 -18520 14796 -17988
rect 14830 -17988 14842 -17944
rect 15800 -17944 15860 -17474
rect 16302 -17732 16362 -17376
rect 16816 -17630 16876 -17286
rect 17836 -17286 17850 -17240
rect 17884 -16768 17898 -16710
rect 18862 -16710 18908 -16698
rect 17884 -17240 17890 -16768
rect 18862 -17230 18868 -16710
rect 17884 -17286 17896 -17240
rect 17114 -17336 17602 -17330
rect 17114 -17370 17126 -17336
rect 17590 -17370 17602 -17336
rect 17114 -17376 17602 -17370
rect 16810 -17690 16816 -17630
rect 16876 -17690 16882 -17630
rect 16300 -17738 16362 -17732
rect 16360 -17798 16362 -17738
rect 16300 -17804 16362 -17798
rect 16812 -17804 16818 -17744
rect 16878 -17804 16884 -17744
rect 16302 -17854 16362 -17804
rect 16096 -17860 16584 -17854
rect 16096 -17894 16108 -17860
rect 16572 -17894 16584 -17860
rect 16096 -17900 16584 -17894
rect 15800 -17988 15814 -17944
rect 14830 -18520 14836 -17988
rect 14790 -18532 14836 -18520
rect 15808 -18520 15814 -17988
rect 15848 -17988 15860 -17944
rect 16818 -17944 16878 -17804
rect 17326 -17854 17386 -17376
rect 17836 -17414 17896 -17286
rect 18854 -17286 18868 -17230
rect 18902 -17230 18908 -16710
rect 19880 -16710 19926 -16698
rect 18902 -17286 18914 -17230
rect 19880 -17242 19886 -16710
rect 18132 -17336 18620 -17330
rect 18132 -17370 18144 -17336
rect 18608 -17370 18620 -17336
rect 18132 -17376 18620 -17370
rect 17830 -17474 17836 -17414
rect 17896 -17474 17902 -17414
rect 17114 -17860 17602 -17854
rect 17114 -17894 17126 -17860
rect 17590 -17894 17602 -17860
rect 17114 -17900 17602 -17894
rect 16818 -17974 16832 -17944
rect 15848 -18520 15854 -17988
rect 16826 -18480 16832 -17974
rect 15808 -18532 15854 -18520
rect 16818 -18520 16832 -18480
rect 16866 -17974 16878 -17944
rect 17836 -17944 17896 -17474
rect 18352 -17854 18412 -17376
rect 18854 -17630 18914 -17286
rect 19870 -17286 19886 -17242
rect 19920 -17242 19926 -16710
rect 20898 -16710 20944 -16698
rect 20898 -17242 20904 -16710
rect 19920 -17286 19930 -17242
rect 19150 -17336 19638 -17330
rect 19150 -17370 19162 -17336
rect 19626 -17370 19638 -17336
rect 19150 -17376 19638 -17370
rect 18848 -17690 18854 -17630
rect 18914 -17690 18920 -17630
rect 19360 -17680 19420 -17376
rect 19870 -17522 19930 -17286
rect 20894 -17286 20904 -17242
rect 20938 -17242 20944 -16710
rect 21916 -16710 21962 -16698
rect 21916 -17236 21922 -16710
rect 20938 -17286 20954 -17242
rect 20168 -17336 20656 -17330
rect 20168 -17370 20180 -17336
rect 20644 -17370 20656 -17336
rect 20168 -17376 20656 -17370
rect 20376 -17520 20436 -17376
rect 19864 -17582 19870 -17522
rect 19930 -17582 19936 -17522
rect 20374 -17526 20436 -17520
rect 20434 -17586 20436 -17526
rect 20374 -17592 20436 -17586
rect 20376 -17680 20436 -17592
rect 20894 -17630 20954 -17286
rect 21910 -17286 21922 -17236
rect 21956 -17236 21962 -16710
rect 22926 -16710 22986 -16544
rect 23028 -16568 23034 -16508
rect 23094 -16568 23100 -16508
rect 23162 -16526 23222 -16238
rect 22926 -16738 22940 -16710
rect 22934 -17228 22940 -16738
rect 21956 -17286 21970 -17236
rect 21186 -17336 21674 -17330
rect 21186 -17370 21198 -17336
rect 21662 -17370 21674 -17336
rect 21186 -17376 21674 -17370
rect 19360 -17740 20436 -17680
rect 20888 -17690 20894 -17630
rect 20954 -17690 20960 -17630
rect 18848 -17804 18854 -17744
rect 18914 -17804 18920 -17744
rect 18132 -17860 18620 -17854
rect 18132 -17894 18144 -17860
rect 18608 -17894 18620 -17860
rect 18132 -17900 18620 -17894
rect 16866 -18480 16872 -17974
rect 17836 -17984 17850 -17944
rect 16866 -18520 16878 -18480
rect 17844 -18486 17850 -17984
rect 14060 -18570 14548 -18564
rect 14060 -18604 14072 -18570
rect 14536 -18604 14548 -18570
rect 14060 -18610 14548 -18604
rect 15078 -18570 15566 -18564
rect 15078 -18604 15090 -18570
rect 15554 -18604 15566 -18570
rect 15078 -18610 15566 -18604
rect 16096 -18570 16584 -18564
rect 16096 -18604 16108 -18570
rect 16572 -18604 16584 -18570
rect 16096 -18610 16584 -18604
rect 14272 -18658 14332 -18610
rect 13760 -18846 13766 -18786
rect 13826 -18846 13832 -18786
rect 14272 -18896 14332 -18718
rect 10202 -19086 10262 -18940
rect 13268 -18956 14332 -18896
rect 15796 -19044 15802 -18984
rect 15862 -19044 15868 -18984
rect 9988 -19092 10476 -19086
rect 9988 -19126 10000 -19092
rect 10464 -19126 10476 -19092
rect 9988 -19132 10476 -19126
rect 11006 -19092 11494 -19086
rect 11006 -19126 11018 -19092
rect 11482 -19126 11494 -19092
rect 11006 -19132 11494 -19126
rect 12024 -19092 12512 -19086
rect 12024 -19126 12036 -19092
rect 12500 -19126 12512 -19092
rect 12024 -19132 12512 -19126
rect 13042 -19092 13530 -19086
rect 13042 -19126 13054 -19092
rect 13518 -19126 13530 -19092
rect 13042 -19132 13530 -19126
rect 14060 -19092 14548 -19086
rect 14060 -19126 14072 -19092
rect 14536 -19126 14548 -19092
rect 14060 -19132 14548 -19126
rect 15078 -19092 15566 -19086
rect 15078 -19126 15090 -19092
rect 15554 -19126 15566 -19092
rect 15078 -19132 15566 -19126
rect 8722 -19752 8728 -19212
rect 9690 -19214 9706 -19176
rect 8682 -19764 8728 -19752
rect 9700 -19752 9706 -19214
rect 9740 -19214 9750 -19176
rect 10718 -19176 10764 -19164
rect 9740 -19752 9746 -19214
rect 10718 -19710 10724 -19176
rect 9700 -19764 9746 -19752
rect 10710 -19752 10724 -19710
rect 10758 -19710 10764 -19176
rect 11736 -19176 11782 -19164
rect 10758 -19752 10770 -19710
rect 11736 -19714 11742 -19176
rect 7952 -19802 8440 -19796
rect 7952 -19836 7964 -19802
rect 8428 -19836 8440 -19802
rect 7952 -19842 8220 -19836
rect 8224 -19842 8440 -19836
rect 8970 -19802 9458 -19796
rect 8970 -19836 8982 -19802
rect 9446 -19836 9458 -19802
rect 8970 -19842 9458 -19836
rect 9988 -19802 10476 -19796
rect 9988 -19836 10000 -19802
rect 10464 -19836 10476 -19802
rect 9988 -19842 10476 -19836
rect 8160 -19898 8220 -19842
rect 9166 -19898 9226 -19842
rect 10210 -19898 10270 -19842
rect 10710 -19892 10770 -19752
rect 11730 -19752 11742 -19714
rect 11776 -19714 11782 -19176
rect 12754 -19176 12800 -19164
rect 11776 -19752 11790 -19714
rect 12754 -19720 12760 -19176
rect 11006 -19802 11494 -19796
rect 11006 -19836 11018 -19802
rect 11482 -19836 11494 -19802
rect 11006 -19842 11494 -19836
rect 8154 -19958 8160 -19898
rect 8220 -19958 8226 -19898
rect 9160 -19958 9166 -19898
rect 9226 -19958 9232 -19898
rect 10204 -19958 10210 -19898
rect 10270 -19958 10276 -19898
rect 10704 -19952 10710 -19892
rect 10770 -19952 10776 -19892
rect 8160 -20320 8220 -19958
rect 9158 -20174 9164 -20114
rect 9224 -20174 9230 -20114
rect 10198 -20174 10204 -20114
rect 10264 -20174 10270 -20114
rect 9164 -20320 9224 -20174
rect 9682 -20278 9688 -20218
rect 9748 -20278 9754 -20218
rect 7952 -20326 8440 -20320
rect 7952 -20360 7964 -20326
rect 8428 -20360 8440 -20326
rect 7952 -20366 8440 -20360
rect 8970 -20326 9458 -20320
rect 8970 -20360 8982 -20326
rect 9446 -20360 9458 -20326
rect 8970 -20366 9458 -20360
rect 7658 -20492 7670 -20410
rect 7664 -20940 7670 -20492
rect 6686 -20986 6700 -20940
rect 5916 -21036 6404 -21030
rect 5916 -21070 5928 -21036
rect 6392 -21070 6404 -21036
rect 5916 -21076 6404 -21070
rect 6106 -21126 6166 -21076
rect 6100 -21186 6106 -21126
rect 6166 -21186 6172 -21126
rect 6640 -21342 6700 -20986
rect 7660 -20986 7670 -20940
rect 7704 -20492 7718 -20410
rect 8682 -20410 8728 -20398
rect 7704 -20940 7710 -20492
rect 7704 -20986 7720 -20940
rect 8682 -20942 8688 -20410
rect 6934 -21036 7422 -21030
rect 6934 -21070 6946 -21036
rect 7410 -21070 7422 -21036
rect 6934 -21076 7422 -21070
rect 7144 -21126 7204 -21076
rect 7138 -21186 7144 -21126
rect 7204 -21186 7210 -21126
rect 6634 -21402 6640 -21342
rect 6700 -21402 6706 -21342
rect 5614 -21500 5620 -21440
rect 5680 -21500 5686 -21440
rect 7144 -21554 7204 -21186
rect 7660 -21440 7720 -20986
rect 8678 -20986 8688 -20942
rect 8722 -20942 8728 -20410
rect 9688 -20410 9748 -20278
rect 10204 -20320 10264 -20174
rect 9988 -20326 10476 -20320
rect 9988 -20360 10000 -20326
rect 10464 -20360 10476 -20326
rect 9988 -20366 10476 -20360
rect 9688 -20474 9706 -20410
rect 8722 -20986 8738 -20942
rect 7952 -21036 8440 -21030
rect 7952 -21070 7964 -21036
rect 8428 -21070 8440 -21036
rect 7952 -21076 8222 -21070
rect 8230 -21076 8440 -21070
rect 8162 -21126 8222 -21076
rect 8678 -21120 8738 -20986
rect 9700 -20986 9706 -20474
rect 9740 -20474 9748 -20410
rect 10710 -20410 10770 -19952
rect 11218 -20114 11278 -19842
rect 11212 -20174 11218 -20114
rect 11278 -20174 11284 -20114
rect 11218 -20320 11278 -20174
rect 11730 -20218 11790 -19752
rect 12746 -19752 12760 -19720
rect 12794 -19720 12800 -19176
rect 13772 -19176 13818 -19164
rect 13772 -19718 13778 -19176
rect 12794 -19752 12806 -19720
rect 12024 -19802 12512 -19796
rect 12024 -19836 12036 -19802
rect 12500 -19836 12512 -19802
rect 12024 -19842 12512 -19836
rect 12226 -20114 12286 -19842
rect 12746 -19892 12806 -19752
rect 13768 -19752 13778 -19718
rect 13812 -19718 13818 -19176
rect 14790 -19176 14836 -19164
rect 13812 -19752 13828 -19718
rect 14790 -19720 14796 -19176
rect 13042 -19802 13530 -19796
rect 13042 -19836 13054 -19802
rect 13518 -19836 13530 -19802
rect 13042 -19842 13530 -19836
rect 12740 -19952 12746 -19892
rect 12806 -19952 12812 -19892
rect 13270 -20114 13330 -19842
rect 12220 -20174 12226 -20114
rect 12286 -20174 12292 -20114
rect 13264 -20174 13270 -20114
rect 13330 -20174 13336 -20114
rect 11724 -20278 11730 -20218
rect 11790 -20278 11796 -20218
rect 11006 -20326 11494 -20320
rect 11006 -20360 11018 -20326
rect 11482 -20360 11494 -20326
rect 11006 -20366 11494 -20360
rect 10710 -20446 10724 -20410
rect 9740 -20986 9746 -20474
rect 10718 -20928 10724 -20446
rect 9700 -20998 9746 -20986
rect 10714 -20986 10724 -20928
rect 10758 -20446 10770 -20410
rect 11730 -20410 11790 -20278
rect 12226 -20320 12286 -20174
rect 13270 -20320 13330 -20174
rect 13768 -20218 13828 -19752
rect 14782 -19752 14796 -19720
rect 14830 -19720 14836 -19176
rect 15802 -19176 15862 -19044
rect 16096 -19092 16584 -19086
rect 16096 -19126 16108 -19092
rect 16572 -19126 16584 -19092
rect 16096 -19132 16584 -19126
rect 14830 -19752 14842 -19720
rect 14060 -19802 14548 -19796
rect 14060 -19836 14072 -19802
rect 14536 -19836 14548 -19802
rect 14060 -19842 14548 -19836
rect 14260 -20114 14320 -19842
rect 14782 -19892 14842 -19752
rect 15802 -19752 15814 -19176
rect 15848 -19752 15862 -19176
rect 16818 -19176 16878 -18520
rect 17838 -18520 17850 -18486
rect 17884 -17984 17896 -17944
rect 18854 -17944 18914 -17804
rect 19360 -17854 19420 -17740
rect 20376 -17854 20436 -17740
rect 20886 -17804 20892 -17744
rect 20952 -17804 20958 -17744
rect 19150 -17860 19638 -17854
rect 19150 -17894 19162 -17860
rect 19626 -17894 19638 -17860
rect 19150 -17900 19638 -17894
rect 20168 -17860 20656 -17854
rect 20168 -17894 20180 -17860
rect 20644 -17894 20656 -17860
rect 20168 -17900 20656 -17894
rect 17884 -18486 17890 -17984
rect 18854 -17986 18868 -17944
rect 17884 -18520 17898 -18486
rect 17114 -18570 17602 -18564
rect 17114 -18604 17126 -18570
rect 17590 -18604 17602 -18570
rect 17114 -18610 17602 -18604
rect 17314 -18880 17374 -18610
rect 17308 -18940 17314 -18880
rect 17374 -18940 17380 -18880
rect 17314 -19086 17374 -18940
rect 17114 -19092 17602 -19086
rect 17114 -19126 17126 -19092
rect 17590 -19126 17602 -19092
rect 17114 -19132 17602 -19126
rect 16818 -19216 16832 -19176
rect 16826 -19720 16832 -19216
rect 15078 -19802 15566 -19796
rect 15078 -19836 15090 -19802
rect 15554 -19836 15566 -19802
rect 15078 -19842 15566 -19836
rect 14776 -19952 14782 -19892
rect 14842 -19952 14848 -19892
rect 15278 -20114 15338 -19842
rect 14254 -20174 14260 -20114
rect 14320 -20174 14326 -20114
rect 15272 -20174 15278 -20114
rect 15338 -20174 15344 -20114
rect 13762 -20278 13768 -20218
rect 13828 -20278 13834 -20218
rect 12024 -20326 12512 -20320
rect 12024 -20360 12036 -20326
rect 12500 -20360 12512 -20326
rect 12024 -20366 12512 -20360
rect 13042 -20326 13530 -20320
rect 13042 -20360 13054 -20326
rect 13518 -20360 13530 -20326
rect 13042 -20366 13530 -20360
rect 10758 -20928 10764 -20446
rect 11730 -20448 11742 -20410
rect 10758 -20986 10774 -20928
rect 8970 -21036 9458 -21030
rect 8970 -21070 8982 -21036
rect 9446 -21070 9458 -21036
rect 8970 -21076 9458 -21070
rect 9988 -21036 10476 -21030
rect 9988 -21070 10000 -21036
rect 10464 -21070 10476 -21036
rect 9988 -21076 10476 -21070
rect 10714 -21120 10774 -20986
rect 11736 -20986 11742 -20448
rect 11776 -20448 11790 -20410
rect 12754 -20410 12800 -20398
rect 11776 -20986 11782 -20448
rect 12754 -20936 12760 -20410
rect 11736 -20998 11782 -20986
rect 12746 -20986 12760 -20936
rect 12794 -20936 12800 -20410
rect 13768 -20410 13828 -20278
rect 14260 -20320 14320 -20174
rect 15802 -20218 15862 -19752
rect 16820 -19752 16832 -19720
rect 16866 -19216 16878 -19176
rect 17838 -19176 17898 -18520
rect 18862 -18520 18868 -17986
rect 18902 -17986 18914 -17944
rect 19880 -17944 19926 -17932
rect 18902 -18520 18908 -17986
rect 19880 -18462 19886 -17944
rect 18862 -18532 18908 -18520
rect 19872 -18520 19886 -18462
rect 19920 -18462 19926 -17944
rect 20892 -17944 20952 -17804
rect 21394 -17854 21454 -17376
rect 21910 -17414 21970 -17286
rect 22928 -17286 22940 -17228
rect 22974 -16738 22986 -16710
rect 22974 -17228 22980 -16738
rect 22974 -17286 22988 -17228
rect 22204 -17336 22692 -17330
rect 22204 -17370 22216 -17336
rect 22680 -17370 22692 -17336
rect 22204 -17376 22692 -17370
rect 22928 -17396 22988 -17286
rect 21904 -17474 21910 -17414
rect 21970 -17474 21976 -17414
rect 22922 -17456 22928 -17396
rect 22988 -17456 22994 -17396
rect 21910 -17692 21970 -17474
rect 21910 -17752 22984 -17692
rect 23034 -17744 23094 -16568
rect 23156 -16586 23162 -16526
rect 23222 -16586 23228 -16526
rect 23528 -17526 23588 -13640
rect 23522 -17586 23528 -17526
rect 23588 -17586 23594 -17526
rect 23272 -17690 23278 -17630
rect 23338 -17690 23344 -17630
rect 21186 -17860 21674 -17854
rect 21186 -17894 21198 -17860
rect 21662 -17894 21674 -17860
rect 21186 -17900 21674 -17894
rect 20892 -17986 20904 -17944
rect 19920 -18520 19932 -18462
rect 18344 -18564 18404 -18562
rect 18132 -18570 18620 -18564
rect 18132 -18604 18144 -18570
rect 18608 -18604 18620 -18570
rect 18132 -18610 18620 -18604
rect 19150 -18570 19638 -18564
rect 19150 -18604 19162 -18570
rect 19626 -18604 19638 -18570
rect 19150 -18610 19638 -18604
rect 18344 -18880 18404 -18610
rect 19366 -18658 19426 -18610
rect 19360 -18718 19366 -18658
rect 19426 -18718 19432 -18658
rect 19498 -18714 19504 -18654
rect 19564 -18714 19570 -18654
rect 19504 -18880 19564 -18714
rect 19872 -18880 19932 -18520
rect 20898 -18520 20904 -17986
rect 20938 -17986 20952 -17944
rect 21910 -17944 21970 -17752
rect 22414 -17854 22474 -17752
rect 22204 -17860 22692 -17854
rect 22204 -17894 22216 -17860
rect 22680 -17894 22692 -17860
rect 22204 -17900 22692 -17894
rect 21910 -17978 21922 -17944
rect 20938 -18520 20944 -17986
rect 21916 -18480 21922 -17978
rect 20898 -18532 20944 -18520
rect 21910 -18520 21922 -18480
rect 21956 -17978 21970 -17944
rect 22924 -17944 22984 -17752
rect 23028 -17804 23034 -17744
rect 23094 -17804 23100 -17744
rect 22924 -17968 22940 -17944
rect 21956 -18480 21962 -17978
rect 21956 -18520 21970 -18480
rect 20168 -18570 20656 -18564
rect 20168 -18604 20180 -18570
rect 20644 -18604 20656 -18570
rect 20168 -18610 20656 -18604
rect 21186 -18570 21674 -18564
rect 21186 -18604 21198 -18570
rect 21662 -18604 21674 -18570
rect 21186 -18610 21674 -18604
rect 21392 -18654 21452 -18610
rect 20380 -18714 20386 -18654
rect 20446 -18714 20452 -18654
rect 21386 -18714 21392 -18654
rect 21452 -18714 21458 -18654
rect 21910 -18658 21970 -18520
rect 22934 -18520 22940 -17968
rect 22974 -17968 22984 -17944
rect 22974 -18520 22980 -17968
rect 22934 -18532 22980 -18520
rect 22204 -18570 22692 -18564
rect 22204 -18604 22216 -18570
rect 22680 -18604 22692 -18570
rect 22204 -18610 22692 -18604
rect 18338 -18940 18344 -18880
rect 18404 -18940 18410 -18880
rect 19498 -18940 19504 -18880
rect 19564 -18940 19570 -18880
rect 19866 -18940 19872 -18880
rect 19932 -18940 19938 -18880
rect 18344 -19086 18404 -18940
rect 19504 -19086 19564 -18940
rect 19872 -18984 19932 -18940
rect 19866 -19044 19872 -18984
rect 19932 -19044 19938 -18984
rect 20386 -19086 20446 -18714
rect 21904 -18718 21910 -18658
rect 21970 -18718 21976 -18658
rect 21904 -18846 21910 -18786
rect 21970 -18846 21976 -18786
rect 20882 -19042 20888 -18982
rect 20948 -19042 20954 -18982
rect 18132 -19092 18620 -19086
rect 18132 -19126 18144 -19092
rect 18608 -19126 18620 -19092
rect 18132 -19132 18620 -19126
rect 19150 -19092 19638 -19086
rect 19150 -19126 19162 -19092
rect 19626 -19126 19638 -19092
rect 19150 -19132 19638 -19126
rect 20168 -19092 20656 -19086
rect 20168 -19126 20180 -19092
rect 20644 -19126 20656 -19092
rect 20168 -19132 20656 -19126
rect 20386 -19134 20446 -19132
rect 16866 -19720 16872 -19216
rect 17838 -19222 17850 -19176
rect 17844 -19708 17850 -19222
rect 16866 -19752 16880 -19720
rect 16096 -19802 16584 -19796
rect 16096 -19836 16108 -19802
rect 16572 -19836 16584 -19802
rect 16096 -19842 16584 -19836
rect 16312 -20114 16372 -19842
rect 16820 -19892 16880 -19752
rect 17836 -19752 17850 -19708
rect 17884 -19222 17898 -19176
rect 18862 -19176 18908 -19164
rect 17884 -19708 17890 -19222
rect 17884 -19752 17896 -19708
rect 18862 -19712 18868 -19176
rect 17114 -19802 17602 -19796
rect 17114 -19836 17126 -19802
rect 17590 -19836 17602 -19802
rect 17114 -19842 17602 -19836
rect 16814 -19952 16820 -19892
rect 16880 -19952 16886 -19892
rect 16806 -20060 16812 -20000
rect 16872 -20060 16878 -20000
rect 16306 -20174 16312 -20114
rect 16372 -20174 16378 -20114
rect 15796 -20278 15802 -20218
rect 15862 -20278 15868 -20218
rect 16308 -20282 16314 -20222
rect 16374 -20282 16380 -20222
rect 16314 -20320 16374 -20282
rect 14060 -20326 14548 -20320
rect 14060 -20360 14072 -20326
rect 14536 -20360 14548 -20326
rect 14060 -20366 14548 -20360
rect 15078 -20326 15566 -20320
rect 15078 -20360 15090 -20326
rect 15554 -20360 15566 -20326
rect 15078 -20366 15566 -20360
rect 16096 -20326 16584 -20320
rect 16096 -20360 16108 -20326
rect 16572 -20360 16584 -20326
rect 16096 -20366 16584 -20360
rect 13768 -20446 13778 -20410
rect 12794 -20986 12806 -20936
rect 11006 -21036 11494 -21030
rect 11006 -21070 11018 -21036
rect 11482 -21070 11494 -21036
rect 11006 -21076 11494 -21070
rect 12024 -21036 12512 -21030
rect 12024 -21070 12036 -21036
rect 12500 -21070 12512 -21036
rect 12024 -21076 12512 -21070
rect 12746 -21120 12806 -20986
rect 13772 -20986 13778 -20446
rect 13812 -20446 13828 -20410
rect 14790 -20410 14836 -20398
rect 13812 -20986 13818 -20446
rect 14790 -20924 14796 -20410
rect 13772 -20998 13818 -20986
rect 14780 -20986 14796 -20924
rect 14830 -20924 14836 -20410
rect 15808 -20410 15854 -20398
rect 14830 -20986 14840 -20924
rect 15808 -20944 15814 -20410
rect 13042 -21036 13530 -21030
rect 13042 -21070 13054 -21036
rect 13518 -21070 13530 -21036
rect 13042 -21076 13530 -21070
rect 14060 -21036 14548 -21030
rect 14060 -21070 14072 -21036
rect 14536 -21070 14548 -21036
rect 14060 -21076 14548 -21070
rect 14780 -21120 14840 -20986
rect 15802 -20986 15814 -20944
rect 15848 -20944 15854 -20410
rect 16812 -20410 16872 -20060
rect 17336 -20222 17396 -19842
rect 17836 -20216 17896 -19752
rect 18856 -19752 18868 -19712
rect 18902 -19712 18908 -19176
rect 19880 -19176 19926 -19164
rect 19880 -19708 19886 -19176
rect 18902 -19752 18916 -19712
rect 18132 -19802 18620 -19796
rect 18132 -19836 18144 -19802
rect 18608 -19836 18620 -19802
rect 18132 -19842 18620 -19836
rect 17330 -20282 17336 -20222
rect 17396 -20282 17402 -20222
rect 17830 -20276 17836 -20216
rect 17896 -20276 17902 -20216
rect 17336 -20320 17396 -20282
rect 17114 -20326 17602 -20320
rect 17114 -20360 17126 -20326
rect 17590 -20360 17602 -20326
rect 17114 -20366 17602 -20360
rect 16812 -20446 16832 -20410
rect 15848 -20986 15862 -20944
rect 15078 -21036 15566 -21030
rect 15078 -21070 15090 -21036
rect 15554 -21070 15566 -21036
rect 15078 -21076 15566 -21070
rect 8156 -21186 8162 -21126
rect 8222 -21186 8228 -21126
rect 8672 -21180 8678 -21120
rect 8738 -21180 8744 -21120
rect 12740 -21180 12746 -21120
rect 12806 -21180 12812 -21120
rect 14774 -21180 14780 -21120
rect 14840 -21180 14846 -21120
rect 7654 -21500 7660 -21440
rect 7720 -21500 7726 -21440
rect 3880 -21560 4368 -21554
rect 3880 -21594 3892 -21560
rect 4356 -21594 4368 -21560
rect 3880 -21600 4368 -21594
rect 4898 -21560 5386 -21554
rect 4898 -21594 4910 -21560
rect 5374 -21594 5386 -21560
rect 4898 -21600 5386 -21594
rect 5916 -21560 6404 -21554
rect 5916 -21594 5928 -21560
rect 6392 -21594 6404 -21560
rect 5916 -21600 6404 -21594
rect 6934 -21560 7422 -21554
rect 6934 -21594 6946 -21560
rect 7410 -21594 7422 -21560
rect 6934 -21600 7422 -21594
rect 3582 -21698 3598 -21644
rect 2614 -22220 2624 -22186
rect 3592 -22190 3598 -21698
rect 2564 -22352 2624 -22220
rect 3588 -22220 3598 -22190
rect 3632 -21698 3642 -21644
rect 4610 -21644 4656 -21632
rect 3632 -22190 3638 -21698
rect 4610 -22174 4616 -21644
rect 3632 -22220 3648 -22190
rect 2862 -22270 3350 -22264
rect 2862 -22304 2874 -22270
rect 3338 -22304 3350 -22270
rect 2862 -22310 3350 -22304
rect 3084 -22352 3144 -22310
rect 3588 -22352 3648 -22220
rect 4602 -22220 4616 -22174
rect 4650 -22174 4656 -21644
rect 5628 -21644 5674 -21632
rect 4650 -22220 4662 -22174
rect 5628 -22190 5634 -21644
rect 3880 -22270 4368 -22264
rect 3880 -22304 3892 -22270
rect 4356 -22304 4368 -22270
rect 3880 -22310 4368 -22304
rect 2564 -22412 3648 -22352
rect 2442 -22522 2448 -22462
rect 2508 -22522 2514 -22462
rect 3588 -22558 3648 -22412
rect 2564 -22618 3648 -22558
rect 2564 -22876 2624 -22618
rect 3076 -22786 3136 -22618
rect 3588 -22678 3648 -22618
rect 3582 -22738 3588 -22678
rect 3648 -22738 3654 -22678
rect 2862 -22792 3350 -22786
rect 2862 -22826 2874 -22792
rect 3338 -22826 3350 -22792
rect 2862 -22832 3350 -22826
rect 2564 -22912 2580 -22876
rect 2574 -23452 2580 -22912
rect 2614 -22912 2624 -22876
rect 3588 -22876 3648 -22738
rect 4080 -22786 4140 -22310
rect 4602 -22364 4662 -22220
rect 5620 -22220 5634 -22190
rect 5668 -22190 5674 -21644
rect 6646 -21644 6692 -21632
rect 6646 -22178 6652 -21644
rect 5668 -22220 5680 -22190
rect 4898 -22270 5386 -22264
rect 4898 -22304 4910 -22270
rect 5374 -22304 5386 -22270
rect 4898 -22310 5386 -22304
rect 4596 -22424 4602 -22364
rect 4662 -22424 4668 -22364
rect 4600 -22618 4606 -22558
rect 4666 -22618 4672 -22558
rect 3880 -22792 4368 -22786
rect 3880 -22826 3892 -22792
rect 4356 -22826 4368 -22792
rect 3880 -22832 4368 -22826
rect 2614 -23452 2620 -22912
rect 3588 -22916 3598 -22876
rect 2574 -23464 2620 -23452
rect 3592 -23452 3598 -22916
rect 3632 -22916 3648 -22876
rect 4606 -22876 4666 -22618
rect 5100 -22622 5160 -22310
rect 5620 -22462 5680 -22220
rect 6638 -22220 6652 -22178
rect 6686 -22178 6692 -21644
rect 7660 -21644 7720 -21500
rect 8162 -21554 8222 -21186
rect 7952 -21560 8440 -21554
rect 7952 -21594 7964 -21560
rect 8428 -21594 8440 -21560
rect 7952 -21600 8440 -21594
rect 7660 -21674 7670 -21644
rect 7664 -22156 7670 -21674
rect 6686 -22220 6698 -22178
rect 5916 -22270 6404 -22264
rect 5916 -22304 5928 -22270
rect 6392 -22304 6404 -22270
rect 5916 -22310 6404 -22304
rect 5614 -22522 5620 -22462
rect 5680 -22522 5686 -22462
rect 6134 -22622 6194 -22310
rect 6638 -22364 6698 -22220
rect 7656 -22220 7670 -22156
rect 7704 -21674 7720 -21644
rect 8678 -21644 8738 -21180
rect 10714 -21186 10774 -21180
rect 11724 -21290 11730 -21230
rect 11790 -21290 11796 -21230
rect 13760 -21290 13766 -21230
rect 13826 -21290 13832 -21230
rect 10706 -21402 10712 -21342
rect 10772 -21402 10778 -21342
rect 9690 -21500 9696 -21440
rect 9756 -21500 9762 -21440
rect 8970 -21560 9458 -21554
rect 8970 -21594 8982 -21560
rect 9446 -21594 9458 -21560
rect 8970 -21600 9458 -21594
rect 7704 -22156 7710 -21674
rect 8678 -21686 8688 -21644
rect 7704 -22220 7716 -22156
rect 8682 -22180 8688 -21686
rect 6934 -22270 7422 -22264
rect 6934 -22304 6946 -22270
rect 7410 -22304 7422 -22270
rect 6934 -22310 7422 -22304
rect 6632 -22424 6638 -22364
rect 6698 -22424 6704 -22364
rect 7144 -22462 7204 -22310
rect 7138 -22522 7144 -22462
rect 7204 -22522 7210 -22462
rect 6636 -22618 6642 -22558
rect 6702 -22618 6708 -22558
rect 5100 -22682 6194 -22622
rect 5100 -22786 5160 -22682
rect 6134 -22786 6194 -22682
rect 4898 -22792 5386 -22786
rect 4898 -22826 4910 -22792
rect 5374 -22826 5386 -22792
rect 4898 -22832 5386 -22826
rect 5916 -22792 6404 -22786
rect 5916 -22826 5928 -22792
rect 6392 -22826 6404 -22792
rect 5916 -22832 6404 -22826
rect 3632 -23452 3638 -22916
rect 4606 -22920 4616 -22876
rect 3592 -23464 3638 -23452
rect 4610 -23452 4616 -22920
rect 4650 -22920 4666 -22876
rect 5628 -22876 5674 -22864
rect 4650 -23452 4656 -22920
rect 5628 -23410 5634 -22876
rect 4610 -23464 4656 -23452
rect 5620 -23452 5634 -23410
rect 5668 -23410 5674 -22876
rect 6642 -22876 6702 -22618
rect 7144 -22786 7204 -22522
rect 7656 -22678 7716 -22220
rect 8676 -22220 8688 -22180
rect 8722 -21686 8738 -21644
rect 9696 -21644 9756 -21500
rect 9988 -21560 10476 -21554
rect 9988 -21594 10000 -21560
rect 10464 -21594 10476 -21560
rect 9988 -21600 10476 -21594
rect 9696 -21680 9706 -21644
rect 8722 -22180 8728 -21686
rect 8722 -22220 8736 -22180
rect 9700 -22186 9706 -21680
rect 7952 -22270 8440 -22264
rect 7952 -22304 7964 -22270
rect 8428 -22304 8440 -22270
rect 7952 -22310 8440 -22304
rect 8166 -22462 8226 -22310
rect 8676 -22364 8736 -22220
rect 9690 -22220 9706 -22186
rect 9740 -21680 9756 -21644
rect 10712 -21644 10772 -21402
rect 11006 -21560 11494 -21554
rect 11006 -21594 11018 -21560
rect 11482 -21594 11494 -21560
rect 11006 -21600 11494 -21594
rect 10712 -21670 10724 -21644
rect 9740 -22186 9746 -21680
rect 10718 -22164 10724 -21670
rect 9740 -22220 9750 -22186
rect 8970 -22270 9458 -22264
rect 8970 -22304 8982 -22270
rect 9446 -22304 9458 -22270
rect 8970 -22310 9458 -22304
rect 8670 -22424 8676 -22364
rect 8736 -22424 8742 -22364
rect 9190 -22456 9250 -22310
rect 7650 -22738 7656 -22678
rect 7716 -22738 7722 -22678
rect 6934 -22792 7422 -22786
rect 6934 -22826 6946 -22792
rect 7410 -22826 7422 -22792
rect 6934 -22832 7422 -22826
rect 6642 -22928 6652 -22876
rect 5668 -23452 5680 -23410
rect 2862 -23502 3350 -23496
rect 2862 -23536 2874 -23502
rect 3338 -23536 3350 -23502
rect 2862 -23542 3350 -23536
rect 3880 -23502 4368 -23496
rect 3880 -23536 3892 -23502
rect 4356 -23536 4368 -23502
rect 3880 -23542 4368 -23536
rect 4898 -23502 5386 -23496
rect 4898 -23536 4910 -23502
rect 5374 -23536 5386 -23502
rect 4898 -23542 5386 -23536
rect 2330 -23654 2336 -23594
rect 2396 -23654 2402 -23594
rect 2224 -23780 2230 -23720
rect 2290 -23780 2296 -23720
rect 2564 -23960 3644 -23900
rect 2564 -24110 2624 -23960
rect 3072 -24020 3132 -23960
rect 2862 -24026 3350 -24020
rect 2862 -24060 2874 -24026
rect 3338 -24060 3350 -24026
rect 2862 -24066 3350 -24060
rect 2564 -24166 2580 -24110
rect 2574 -24592 2580 -24166
rect 2614 -24166 2624 -24110
rect 3584 -24110 3644 -23960
rect 4082 -24020 4142 -23542
rect 5620 -23720 5680 -23452
rect 6646 -23452 6652 -22928
rect 6686 -22928 6702 -22876
rect 7656 -22876 7716 -22738
rect 8166 -22786 8226 -22522
rect 9188 -22462 9250 -22456
rect 9248 -22522 9250 -22462
rect 9188 -22528 9250 -22522
rect 8664 -22618 8670 -22558
rect 8730 -22618 8736 -22558
rect 7952 -22792 8440 -22786
rect 7952 -22826 7964 -22792
rect 8428 -22826 8440 -22792
rect 7952 -22832 8440 -22826
rect 7656 -22916 7670 -22876
rect 6686 -23452 6692 -22928
rect 7664 -23398 7670 -22916
rect 6646 -23464 6692 -23452
rect 7658 -23452 7670 -23398
rect 7704 -22916 7716 -22876
rect 8670 -22876 8730 -22618
rect 9190 -22786 9250 -22528
rect 9690 -22678 9750 -22220
rect 10708 -22220 10724 -22164
rect 10758 -21670 10772 -21644
rect 11730 -21644 11790 -21290
rect 12024 -21560 12512 -21554
rect 12024 -21594 12036 -21560
rect 12500 -21594 12512 -21560
rect 12024 -21600 12512 -21594
rect 13042 -21560 13530 -21554
rect 13042 -21594 13054 -21560
rect 13518 -21594 13530 -21560
rect 13042 -21600 13530 -21594
rect 10758 -22164 10764 -21670
rect 11730 -21676 11742 -21644
rect 10758 -22220 10768 -22164
rect 9988 -22270 10476 -22264
rect 9988 -22304 10000 -22270
rect 10464 -22304 10476 -22270
rect 9988 -22310 10252 -22304
rect 10264 -22310 10476 -22304
rect 10192 -22462 10252 -22310
rect 10538 -22344 10598 -22338
rect 10708 -22344 10768 -22220
rect 11736 -22220 11742 -21676
rect 11776 -21676 11790 -21644
rect 12754 -21644 12800 -21632
rect 11776 -22220 11782 -21676
rect 12754 -22150 12760 -21644
rect 11736 -22232 11782 -22220
rect 12750 -22220 12760 -22150
rect 12794 -22150 12800 -21644
rect 13766 -21644 13826 -21290
rect 15308 -21328 15368 -21076
rect 15802 -21118 15862 -20986
rect 16826 -20986 16832 -20446
rect 16866 -20986 16872 -20410
rect 17836 -20410 17896 -20276
rect 18314 -20320 18374 -19842
rect 18856 -19892 18916 -19752
rect 19870 -19752 19886 -19708
rect 19920 -19708 19926 -19176
rect 20888 -19176 20948 -19042
rect 21186 -19092 21674 -19086
rect 21186 -19126 21198 -19092
rect 21662 -19126 21674 -19092
rect 21186 -19132 21674 -19126
rect 20888 -19226 20904 -19176
rect 19920 -19752 19930 -19708
rect 20898 -19724 20904 -19226
rect 19150 -19802 19638 -19796
rect 19150 -19836 19162 -19802
rect 19626 -19836 19638 -19802
rect 19150 -19842 19638 -19836
rect 18850 -19952 18856 -19892
rect 18916 -19952 18922 -19892
rect 18846 -20060 18852 -20000
rect 18912 -20060 18918 -20000
rect 18132 -20326 18620 -20320
rect 18132 -20360 18144 -20326
rect 18608 -20360 18620 -20326
rect 18132 -20366 18620 -20360
rect 17836 -20504 17850 -20410
rect 17844 -20944 17850 -20504
rect 16826 -20998 16872 -20986
rect 17836 -20986 17850 -20944
rect 17884 -20504 17896 -20410
rect 18852 -20410 18912 -20060
rect 19338 -20174 19344 -20114
rect 19404 -20174 19410 -20114
rect 19344 -20320 19404 -20174
rect 19870 -20216 19930 -19752
rect 20894 -19752 20904 -19724
rect 20938 -19226 20948 -19176
rect 21910 -19176 21970 -18846
rect 22204 -19092 22692 -19086
rect 22204 -19126 22216 -19092
rect 22680 -19126 22692 -19092
rect 22204 -19132 22692 -19126
rect 20938 -19724 20944 -19226
rect 21910 -19228 21922 -19176
rect 21916 -19724 21922 -19228
rect 20938 -19752 20954 -19724
rect 20168 -19802 20656 -19796
rect 20168 -19836 20180 -19802
rect 20644 -19836 20656 -19802
rect 20168 -19842 20656 -19836
rect 20894 -19892 20954 -19752
rect 21910 -19752 21922 -19724
rect 21956 -19228 21970 -19176
rect 22934 -19176 22980 -19164
rect 21956 -19724 21962 -19228
rect 22934 -19718 22940 -19176
rect 21956 -19752 21970 -19724
rect 21186 -19802 21674 -19796
rect 21186 -19836 21198 -19802
rect 21662 -19836 21674 -19802
rect 21186 -19842 21674 -19836
rect 20888 -19952 20894 -19892
rect 20954 -19952 20960 -19892
rect 20884 -20060 20890 -20000
rect 20950 -20060 20956 -20000
rect 20376 -20174 20382 -20114
rect 20442 -20174 20448 -20114
rect 19864 -20276 19870 -20216
rect 19930 -20276 19936 -20216
rect 20382 -20320 20442 -20174
rect 19150 -20326 19638 -20320
rect 19150 -20360 19162 -20326
rect 19626 -20360 19638 -20326
rect 19150 -20366 19638 -20360
rect 20168 -20326 20656 -20320
rect 20168 -20360 20180 -20326
rect 20644 -20360 20656 -20326
rect 20168 -20366 20656 -20360
rect 18852 -20476 18868 -20410
rect 17884 -20944 17890 -20504
rect 17884 -20986 17896 -20944
rect 16096 -21036 16584 -21030
rect 16096 -21070 16108 -21036
rect 16572 -21070 16584 -21036
rect 16096 -21076 16584 -21070
rect 17114 -21036 17602 -21030
rect 17114 -21070 17126 -21036
rect 17590 -21070 17602 -21036
rect 17114 -21076 17602 -21070
rect 15796 -21178 15802 -21118
rect 15862 -21178 15868 -21118
rect 16150 -21178 16156 -21118
rect 16216 -21178 16222 -21118
rect 15792 -21290 15798 -21230
rect 15858 -21290 15864 -21230
rect 15302 -21388 15308 -21328
rect 15368 -21388 15374 -21328
rect 14060 -21560 14548 -21554
rect 14060 -21594 14072 -21560
rect 14536 -21594 14548 -21560
rect 14060 -21600 14548 -21594
rect 15078 -21560 15566 -21554
rect 15078 -21594 15090 -21560
rect 15554 -21594 15566 -21560
rect 15078 -21600 15566 -21594
rect 13766 -21682 13778 -21644
rect 12794 -22220 12810 -22150
rect 11006 -22270 11494 -22264
rect 11006 -22304 11018 -22270
rect 11482 -22304 11494 -22270
rect 11006 -22310 11494 -22304
rect 12024 -22270 12512 -22264
rect 12024 -22304 12036 -22270
rect 12500 -22304 12512 -22270
rect 12024 -22310 12512 -22304
rect 10702 -22404 10708 -22344
rect 10768 -22404 10774 -22344
rect 10186 -22522 10192 -22462
rect 10252 -22522 10258 -22462
rect 9684 -22738 9690 -22678
rect 9750 -22738 9756 -22678
rect 8970 -22792 9458 -22786
rect 8970 -22826 8982 -22792
rect 9446 -22826 9458 -22792
rect 8970 -22832 9458 -22826
rect 7704 -23398 7710 -22916
rect 8670 -22936 8688 -22876
rect 7704 -23452 7718 -23398
rect 5916 -23502 6404 -23496
rect 5916 -23536 5928 -23502
rect 6392 -23536 6404 -23502
rect 5916 -23542 6256 -23536
rect 6316 -23542 6404 -23536
rect 6934 -23502 7422 -23496
rect 6934 -23536 6946 -23502
rect 7410 -23536 7422 -23502
rect 6934 -23542 7422 -23536
rect 6140 -23708 6200 -23542
rect 5614 -23780 5620 -23720
rect 5680 -23780 5686 -23720
rect 6134 -23768 6140 -23708
rect 6200 -23768 6206 -23708
rect 4596 -23882 4602 -23822
rect 4662 -23882 4668 -23822
rect 6632 -23882 6638 -23822
rect 6698 -23882 6704 -23822
rect 3880 -24026 4368 -24020
rect 3880 -24060 3892 -24026
rect 4356 -24060 4368 -24026
rect 3880 -24066 4368 -24060
rect 2614 -24592 2620 -24166
rect 3584 -24686 3598 -24110
rect 3632 -24686 3644 -24110
rect 4602 -24110 4662 -23882
rect 5614 -23986 5620 -23926
rect 5680 -23986 5686 -23926
rect 4898 -24026 5386 -24020
rect 4898 -24060 4910 -24026
rect 5374 -24060 5386 -24026
rect 4898 -24066 5386 -24060
rect 4602 -24170 4616 -24110
rect 4610 -24592 4616 -24170
rect 2442 -24884 2448 -24824
rect 2508 -24884 2514 -24824
rect 2114 -24988 2120 -24928
rect 2180 -24988 2186 -24928
rect 2448 -25154 2508 -24884
rect 3584 -24928 3644 -24686
rect 4604 -24686 4616 -24650
rect 4650 -24170 4662 -24110
rect 5620 -24110 5680 -23986
rect 5916 -24026 6140 -24020
rect 6200 -24026 6256 -24020
rect 6316 -24026 6404 -24020
rect 5916 -24060 5928 -24026
rect 6392 -24060 6404 -24026
rect 5916 -24066 6404 -24060
rect 5620 -24164 5634 -24110
rect 4650 -24592 4656 -24170
rect 5628 -24592 5634 -24164
rect 4650 -24686 4664 -24650
rect 3578 -24988 3584 -24928
rect 3644 -24988 3650 -24928
rect 4092 -25034 4152 -24770
rect 4086 -25094 4092 -25034
rect 4152 -25094 4158 -25034
rect 2448 -25214 3648 -25154
rect 1064 -26048 1070 -25988
rect 1130 -26048 1136 -25988
rect 2448 -26066 2508 -25214
rect 2568 -25414 2628 -25214
rect 3054 -25298 3114 -25214
rect 3588 -25418 3648 -25214
rect 4092 -25288 4152 -25094
rect 4604 -25144 4664 -24686
rect 5618 -24686 5634 -24646
rect 5668 -24164 5680 -24110
rect 6638 -24110 6698 -23882
rect 7140 -24020 7200 -23542
rect 7658 -23822 7718 -23452
rect 8682 -23452 8688 -22936
rect 8722 -22936 8730 -22876
rect 9690 -22876 9750 -22738
rect 10192 -22786 10252 -22522
rect 10538 -22558 10598 -22404
rect 10532 -22618 10538 -22558
rect 10598 -22618 10604 -22558
rect 10708 -22612 10714 -22552
rect 10774 -22612 10780 -22552
rect 9988 -22792 10252 -22786
rect 10264 -22792 10476 -22786
rect 9988 -22826 10000 -22792
rect 10464 -22826 10476 -22792
rect 9988 -22832 10476 -22826
rect 9690 -22916 9706 -22876
rect 8722 -23452 8728 -22936
rect 9700 -23386 9706 -22916
rect 8682 -23464 8728 -23452
rect 9694 -23452 9706 -23386
rect 9740 -22916 9750 -22876
rect 10714 -22876 10774 -22612
rect 11230 -22614 11290 -22310
rect 12244 -22450 12304 -22310
rect 12750 -22344 12810 -22220
rect 13772 -22220 13778 -21682
rect 13812 -21682 13826 -21644
rect 14790 -21644 14836 -21632
rect 13812 -22220 13818 -21682
rect 14790 -22150 14796 -21644
rect 13772 -22232 13818 -22220
rect 14782 -22220 14796 -22150
rect 14830 -22150 14836 -21644
rect 15798 -21644 15858 -21290
rect 16156 -21436 16216 -21178
rect 16346 -21328 16406 -21076
rect 17322 -21328 17382 -21076
rect 16340 -21388 16346 -21328
rect 16406 -21388 16412 -21328
rect 17316 -21388 17322 -21328
rect 17382 -21388 17388 -21328
rect 17836 -21440 17896 -20986
rect 18862 -20986 18868 -20476
rect 18902 -20476 18912 -20410
rect 19880 -20410 19926 -20398
rect 18902 -20986 18908 -20476
rect 19880 -20942 19886 -20410
rect 18862 -20998 18908 -20986
rect 19874 -20986 19886 -20942
rect 19920 -20942 19926 -20410
rect 20890 -20410 20950 -20060
rect 21408 -20114 21468 -19842
rect 21910 -19934 21970 -19752
rect 22924 -19752 22940 -19718
rect 22974 -19718 22980 -19176
rect 22974 -19752 22984 -19718
rect 22204 -19802 22692 -19796
rect 22204 -19836 22216 -19802
rect 22680 -19836 22692 -19802
rect 22204 -19842 22692 -19836
rect 22418 -19934 22478 -19842
rect 22924 -19934 22984 -19752
rect 21910 -19994 22984 -19934
rect 21402 -20174 21408 -20114
rect 21468 -20174 21474 -20114
rect 21906 -20276 21912 -20216
rect 21972 -20276 21978 -20216
rect 21186 -20326 21674 -20320
rect 21186 -20360 21198 -20326
rect 21662 -20360 21674 -20326
rect 21186 -20366 21674 -20360
rect 20890 -20462 20904 -20410
rect 20898 -20936 20904 -20462
rect 19920 -20986 19934 -20942
rect 18132 -21036 18620 -21030
rect 18132 -21070 18144 -21036
rect 18608 -21070 18620 -21036
rect 18132 -21076 18620 -21070
rect 19150 -21036 19638 -21030
rect 19150 -21070 19162 -21036
rect 19626 -21070 19638 -21036
rect 19150 -21076 19638 -21070
rect 18338 -21328 18398 -21076
rect 19874 -21118 19934 -20986
rect 20892 -20986 20904 -20936
rect 20938 -20462 20950 -20410
rect 21912 -20410 21972 -20276
rect 22204 -20326 22692 -20320
rect 22204 -20360 22216 -20326
rect 22680 -20360 22692 -20326
rect 22204 -20366 22692 -20360
rect 21912 -20444 21922 -20410
rect 20938 -20936 20944 -20462
rect 20938 -20986 20952 -20936
rect 21916 -20942 21922 -20444
rect 20168 -21036 20656 -21030
rect 20168 -21070 20180 -21036
rect 20644 -21070 20656 -21036
rect 20168 -21076 20656 -21070
rect 19868 -21178 19874 -21118
rect 19934 -21178 19940 -21118
rect 18332 -21388 18338 -21328
rect 18398 -21388 18404 -21328
rect 20358 -21388 20364 -21328
rect 20424 -21388 20430 -21328
rect 16156 -21502 16216 -21496
rect 17830 -21500 17836 -21440
rect 17896 -21500 17902 -21440
rect 19866 -21500 19872 -21440
rect 19932 -21500 19938 -21440
rect 16096 -21560 16584 -21554
rect 16096 -21594 16108 -21560
rect 16572 -21594 16584 -21560
rect 16096 -21600 16584 -21594
rect 17114 -21560 17602 -21554
rect 17114 -21594 17126 -21560
rect 17590 -21594 17602 -21560
rect 17114 -21600 17602 -21594
rect 15798 -21686 15814 -21644
rect 14830 -22220 14842 -22150
rect 13042 -22270 13530 -22264
rect 13042 -22304 13054 -22270
rect 13518 -22304 13530 -22270
rect 13042 -22310 13530 -22304
rect 14060 -22270 14548 -22264
rect 14060 -22304 14072 -22270
rect 14536 -22304 14548 -22270
rect 14060 -22310 14548 -22304
rect 12744 -22404 12750 -22344
rect 12810 -22404 12816 -22344
rect 13266 -22450 13326 -22310
rect 14280 -22450 14340 -22310
rect 14782 -22344 14842 -22220
rect 15808 -22220 15814 -21686
rect 15848 -21686 15858 -21644
rect 16826 -21644 16872 -21632
rect 15848 -22220 15854 -21686
rect 16826 -22184 16832 -21644
rect 15808 -22232 15854 -22220
rect 16822 -22220 16832 -22184
rect 16866 -22184 16872 -21644
rect 17836 -21644 17896 -21500
rect 18132 -21560 18620 -21554
rect 18132 -21594 18144 -21560
rect 18608 -21594 18620 -21560
rect 18132 -21600 18620 -21594
rect 19150 -21560 19638 -21554
rect 19150 -21594 19162 -21560
rect 19626 -21594 19638 -21560
rect 19150 -21600 19638 -21594
rect 17836 -21682 17850 -21644
rect 17844 -22168 17850 -21682
rect 16866 -22220 16882 -22184
rect 15078 -22270 15566 -22264
rect 15078 -22304 15090 -22270
rect 15554 -22304 15566 -22270
rect 15078 -22310 15566 -22304
rect 16096 -22270 16584 -22264
rect 16096 -22304 16108 -22270
rect 16572 -22304 16584 -22270
rect 16096 -22310 16584 -22304
rect 14776 -22404 14782 -22344
rect 14842 -22404 14848 -22344
rect 15282 -22350 15342 -22310
rect 16308 -22350 16368 -22310
rect 16822 -22344 16882 -22220
rect 17840 -22220 17850 -22168
rect 17884 -21682 17896 -21644
rect 18862 -21644 18908 -21632
rect 17884 -22168 17890 -21682
rect 17884 -22220 17900 -22168
rect 18862 -22176 18868 -21644
rect 17114 -22270 17602 -22264
rect 17114 -22304 17126 -22270
rect 17590 -22304 17602 -22270
rect 17114 -22310 17602 -22304
rect 15282 -22410 16368 -22350
rect 16816 -22404 16822 -22344
rect 16882 -22404 16888 -22344
rect 15282 -22450 15342 -22410
rect 12244 -22510 15342 -22450
rect 15794 -22502 15800 -22442
rect 15860 -22502 15866 -22442
rect 12244 -22614 12304 -22510
rect 12736 -22612 12742 -22552
rect 12802 -22612 12808 -22552
rect 11230 -22674 12304 -22614
rect 11230 -22786 11290 -22674
rect 12244 -22786 12304 -22674
rect 11006 -22792 11494 -22786
rect 11006 -22826 11018 -22792
rect 11482 -22826 11494 -22792
rect 11006 -22832 11494 -22826
rect 12024 -22792 12512 -22786
rect 12024 -22826 12036 -22792
rect 12500 -22826 12512 -22792
rect 12024 -22832 12512 -22826
rect 9740 -23386 9746 -22916
rect 10714 -22920 10724 -22876
rect 9740 -23452 9754 -23386
rect 10718 -23394 10724 -22920
rect 7952 -23502 8440 -23496
rect 7952 -23536 7964 -23502
rect 8428 -23536 8440 -23502
rect 7952 -23542 8440 -23536
rect 8970 -23502 9458 -23496
rect 8970 -23536 8982 -23502
rect 9446 -23536 9458 -23502
rect 8970 -23542 9458 -23536
rect 7652 -23882 7658 -23822
rect 7718 -23882 7724 -23822
rect 8162 -24020 8222 -23542
rect 8668 -23882 8674 -23822
rect 8734 -23882 8740 -23822
rect 6934 -24026 7422 -24020
rect 6934 -24060 6946 -24026
rect 7410 -24060 7422 -24026
rect 6934 -24066 7422 -24060
rect 7952 -24026 8440 -24020
rect 7952 -24060 7964 -24026
rect 8428 -24060 8440 -24026
rect 7952 -24066 8440 -24060
rect 6638 -24160 6652 -24110
rect 5668 -24592 5674 -24164
rect 6646 -24592 6652 -24160
rect 5668 -24686 5678 -24646
rect 5112 -25034 5172 -24770
rect 5618 -24824 5678 -24686
rect 6640 -24686 6652 -24662
rect 6686 -24160 6698 -24110
rect 7664 -24110 7710 -24098
rect 6686 -24592 6692 -24160
rect 7664 -24592 7670 -24110
rect 6686 -24686 6700 -24662
rect 5612 -24884 5618 -24824
rect 5678 -24884 5684 -24824
rect 5618 -24988 5624 -24928
rect 5684 -24988 5690 -24928
rect 5106 -25094 5112 -25034
rect 5172 -25094 5178 -25034
rect 4598 -25204 4604 -25144
rect 4664 -25204 4670 -25144
rect 3584 -26066 3644 -25870
rect 2442 -26126 2448 -26066
rect 2508 -26126 2514 -26066
rect 3578 -26126 3584 -26066
rect 3644 -26126 3650 -26066
rect 4096 -26174 4156 -25970
rect 4090 -26234 4096 -26174
rect 4156 -26234 4162 -26174
rect 4604 -26430 4664 -25204
rect 5112 -25284 5172 -25094
rect 5624 -25356 5684 -24988
rect 6136 -25034 6196 -24770
rect 6130 -25094 6136 -25034
rect 6196 -25094 6202 -25034
rect 6136 -25290 6196 -25094
rect 6640 -25144 6700 -24686
rect 7654 -24686 7670 -24672
rect 7704 -24592 7710 -24110
rect 8674 -24110 8734 -23882
rect 9174 -24020 9234 -23542
rect 9694 -23822 9754 -23452
rect 10706 -23452 10724 -23394
rect 10758 -22920 10774 -22876
rect 11736 -22876 11782 -22864
rect 10758 -23394 10764 -22920
rect 10758 -23452 10766 -23394
rect 11736 -23400 11742 -22876
rect 9988 -23502 10476 -23496
rect 9988 -23536 10000 -23502
rect 10464 -23536 10476 -23502
rect 9988 -23542 10476 -23536
rect 9688 -23882 9694 -23822
rect 9754 -23882 9760 -23822
rect 10204 -24020 10264 -23542
rect 10706 -23654 10766 -23452
rect 11724 -23452 11742 -23400
rect 11776 -23400 11782 -22876
rect 12742 -22876 12802 -22612
rect 13266 -22786 13326 -22510
rect 14280 -22786 14340 -22510
rect 14780 -22612 14786 -22552
rect 14846 -22612 14852 -22552
rect 13042 -22792 13530 -22786
rect 13042 -22826 13054 -22792
rect 13518 -22826 13530 -22792
rect 13042 -22832 13530 -22826
rect 14060 -22792 14548 -22786
rect 14060 -22826 14072 -22792
rect 14536 -22826 14548 -22792
rect 14060 -22832 14548 -22826
rect 12742 -22920 12760 -22876
rect 11776 -23452 11784 -23400
rect 11006 -23502 11494 -23496
rect 11006 -23536 11018 -23502
rect 11482 -23536 11494 -23502
rect 11006 -23542 11494 -23536
rect 10556 -23714 10766 -23654
rect 11220 -23708 11280 -23542
rect 11724 -23594 11784 -23452
rect 12754 -23452 12760 -22920
rect 12794 -22920 12802 -22876
rect 13772 -22876 13818 -22864
rect 12794 -23452 12800 -22920
rect 13772 -23400 13778 -22876
rect 12754 -23464 12800 -23452
rect 13766 -23452 13778 -23400
rect 13812 -23400 13818 -22876
rect 14786 -22876 14846 -22612
rect 15282 -22786 15342 -22510
rect 15078 -22792 15566 -22786
rect 15078 -22826 15090 -22792
rect 15554 -22826 15566 -22792
rect 15078 -22832 15566 -22826
rect 14786 -22924 14796 -22876
rect 13812 -23452 13826 -23400
rect 12024 -23502 12512 -23496
rect 12024 -23536 12036 -23502
rect 12500 -23536 12512 -23502
rect 12024 -23542 12512 -23536
rect 13042 -23502 13530 -23496
rect 13042 -23536 13054 -23502
rect 13518 -23536 13530 -23502
rect 13042 -23542 13530 -23536
rect 13766 -23594 13826 -23452
rect 14790 -23452 14796 -22924
rect 14830 -22924 14846 -22876
rect 15800 -22876 15860 -22502
rect 16308 -22786 16368 -22410
rect 16808 -22612 16814 -22552
rect 16874 -22612 16880 -22552
rect 16096 -22792 16584 -22786
rect 16096 -22826 16108 -22792
rect 16572 -22826 16584 -22792
rect 16096 -22832 16584 -22826
rect 15800 -22912 15814 -22876
rect 14830 -23452 14836 -22924
rect 15808 -23408 15814 -22912
rect 14790 -23464 14836 -23452
rect 15802 -23452 15814 -23408
rect 15848 -22912 15860 -22876
rect 16814 -22876 16874 -22612
rect 17328 -22786 17388 -22310
rect 17840 -22678 17900 -22220
rect 18852 -22220 18868 -22176
rect 18902 -22176 18908 -21644
rect 19872 -21644 19932 -21500
rect 20364 -21554 20424 -21388
rect 20168 -21560 20656 -21554
rect 20168 -21594 20180 -21560
rect 20644 -21594 20656 -21560
rect 20168 -21600 20656 -21594
rect 19872 -21702 19886 -21644
rect 18902 -22220 18912 -22176
rect 19880 -22180 19886 -21702
rect 18132 -22270 18620 -22264
rect 18132 -22304 18144 -22270
rect 18608 -22304 18620 -22270
rect 18132 -22310 18620 -22304
rect 17834 -22738 17840 -22678
rect 17900 -22738 17906 -22678
rect 17114 -22792 17602 -22786
rect 17114 -22826 17126 -22792
rect 17590 -22826 17602 -22792
rect 17114 -22832 17602 -22826
rect 15848 -23408 15854 -22912
rect 16814 -22924 16832 -22876
rect 15848 -23452 15862 -23408
rect 16826 -23412 16832 -22924
rect 14060 -23502 14548 -23496
rect 14060 -23536 14072 -23502
rect 14536 -23536 14548 -23502
rect 14060 -23542 14548 -23536
rect 15078 -23502 15566 -23496
rect 15078 -23536 15090 -23502
rect 15554 -23536 15566 -23502
rect 15078 -23542 15566 -23536
rect 15802 -23594 15862 -23452
rect 16816 -23452 16832 -23412
rect 16866 -22924 16874 -22876
rect 17840 -22876 17900 -22738
rect 18344 -22786 18404 -22310
rect 18852 -22552 18912 -22220
rect 19870 -22220 19886 -22180
rect 19920 -21702 19932 -21644
rect 20892 -21644 20952 -20986
rect 21908 -20986 21922 -20942
rect 21956 -20444 21972 -20410
rect 22934 -20410 22980 -20398
rect 21956 -20942 21962 -20444
rect 21956 -20986 21968 -20942
rect 22934 -20956 22940 -20410
rect 21186 -21036 21674 -21030
rect 21186 -21070 21198 -21036
rect 21662 -21070 21674 -21036
rect 21186 -21076 21674 -21070
rect 21394 -21328 21454 -21076
rect 21908 -21168 21968 -20986
rect 22924 -20986 22940 -20956
rect 22974 -20956 22980 -20410
rect 22974 -20986 22984 -20956
rect 22204 -21036 22692 -21030
rect 22204 -21070 22216 -21036
rect 22680 -21070 22692 -21036
rect 22204 -21076 22692 -21070
rect 22414 -21168 22474 -21076
rect 22924 -21168 22984 -20986
rect 21908 -21228 22984 -21168
rect 21388 -21388 21394 -21328
rect 21454 -21388 21460 -21328
rect 21908 -21440 21968 -21228
rect 21902 -21500 21908 -21440
rect 21968 -21500 21974 -21440
rect 21186 -21560 21674 -21554
rect 21186 -21594 21198 -21560
rect 21662 -21594 21674 -21560
rect 21186 -21600 21674 -21594
rect 22204 -21560 22692 -21554
rect 22204 -21594 22216 -21560
rect 22680 -21594 22692 -21560
rect 22204 -21600 22692 -21594
rect 20892 -21686 20904 -21644
rect 19920 -22180 19926 -21702
rect 20898 -22166 20904 -21686
rect 19920 -22220 19930 -22180
rect 19150 -22270 19638 -22264
rect 19150 -22304 19162 -22270
rect 19626 -22304 19638 -22270
rect 19150 -22310 19638 -22304
rect 18846 -22612 18852 -22552
rect 18912 -22612 18918 -22552
rect 19378 -22786 19438 -22310
rect 19870 -22678 19930 -22220
rect 20892 -22220 20904 -22166
rect 20938 -21686 20952 -21644
rect 21916 -21644 21962 -21632
rect 20938 -22166 20944 -21686
rect 20938 -22220 20952 -22166
rect 21916 -22174 21922 -21644
rect 20168 -22270 20656 -22264
rect 20168 -22304 20180 -22270
rect 20644 -22304 20656 -22270
rect 20168 -22310 20656 -22304
rect 20396 -22676 20456 -22310
rect 20892 -22552 20952 -22220
rect 21906 -22220 21922 -22174
rect 21956 -22174 21962 -21644
rect 22934 -21644 22980 -21632
rect 21956 -22220 21966 -22174
rect 22934 -22192 22940 -21644
rect 21186 -22270 21674 -22264
rect 21186 -22304 21198 -22270
rect 21662 -22304 21674 -22270
rect 21186 -22310 21674 -22304
rect 21410 -22548 21470 -22310
rect 21906 -22346 21966 -22220
rect 22926 -22220 22940 -22192
rect 22974 -22192 22980 -21644
rect 22974 -22220 22986 -22192
rect 22204 -22270 22692 -22264
rect 22204 -22304 22216 -22270
rect 22680 -22304 22692 -22270
rect 22204 -22310 22692 -22304
rect 22412 -22344 22472 -22310
rect 22926 -22344 22986 -22220
rect 22412 -22346 22986 -22344
rect 21906 -22406 22986 -22346
rect 21906 -22442 21966 -22406
rect 21900 -22502 21906 -22442
rect 21966 -22502 21972 -22442
rect 20886 -22612 20892 -22552
rect 20952 -22612 20958 -22552
rect 21404 -22608 21410 -22548
rect 21470 -22608 21476 -22548
rect 22916 -22608 22922 -22548
rect 22982 -22608 22988 -22548
rect 19864 -22738 19870 -22678
rect 19930 -22738 19936 -22678
rect 18132 -22792 18620 -22786
rect 18132 -22826 18144 -22792
rect 18608 -22826 18620 -22792
rect 18132 -22832 18620 -22826
rect 19150 -22792 19638 -22786
rect 19150 -22826 19162 -22792
rect 19626 -22826 19638 -22792
rect 19150 -22832 19638 -22826
rect 17840 -22922 17850 -22876
rect 16866 -23412 16872 -22924
rect 17844 -23392 17850 -22922
rect 16866 -23452 16876 -23412
rect 16096 -23502 16584 -23496
rect 16096 -23536 16108 -23502
rect 16572 -23536 16584 -23502
rect 16096 -23542 16584 -23536
rect 11718 -23654 11724 -23594
rect 11784 -23654 11790 -23594
rect 13760 -23654 13766 -23594
rect 13826 -23654 13832 -23594
rect 15796 -23654 15802 -23594
rect 15862 -23654 15868 -23594
rect 16308 -23704 16368 -23542
rect 16816 -23602 16876 -23452
rect 17838 -23452 17850 -23392
rect 17884 -22922 17900 -22876
rect 18862 -22876 18908 -22864
rect 17884 -23392 17890 -22922
rect 17884 -23452 17898 -23392
rect 18862 -23408 18868 -22876
rect 17114 -23502 17602 -23496
rect 17114 -23536 17126 -23502
rect 17590 -23536 17602 -23502
rect 17114 -23542 17602 -23536
rect 16816 -23662 17022 -23602
rect 10556 -23926 10616 -23714
rect 11214 -23768 11220 -23708
rect 11280 -23768 11286 -23708
rect 16302 -23764 16308 -23704
rect 16368 -23764 16374 -23704
rect 10706 -23882 10712 -23822
rect 10772 -23882 10778 -23822
rect 12736 -23882 12742 -23822
rect 12802 -23882 12808 -23822
rect 14774 -23882 14780 -23822
rect 14840 -23882 14846 -23822
rect 16810 -23882 16816 -23822
rect 16876 -23882 16882 -23822
rect 10550 -23986 10556 -23926
rect 10616 -23986 10622 -23926
rect 8970 -24026 9458 -24020
rect 8970 -24060 8982 -24026
rect 9446 -24060 9458 -24026
rect 8970 -24066 9458 -24060
rect 9988 -24026 10476 -24020
rect 9988 -24060 10000 -24026
rect 10464 -24060 10476 -24026
rect 9988 -24066 10476 -24060
rect 8674 -24592 8688 -24110
rect 7704 -24686 7714 -24672
rect 7154 -25034 7214 -24770
rect 7654 -24928 7714 -24686
rect 8678 -24686 8688 -24666
rect 8722 -24592 8734 -24110
rect 9700 -24110 9746 -24098
rect 9700 -24592 9706 -24110
rect 8722 -24686 8738 -24666
rect 7648 -24988 7654 -24928
rect 7714 -24988 7720 -24928
rect 8168 -25034 8228 -24770
rect 7148 -25094 7154 -25034
rect 7214 -25094 7220 -25034
rect 8162 -25094 8168 -25034
rect 8228 -25094 8234 -25034
rect 6634 -25204 6640 -25144
rect 6700 -25204 6706 -25144
rect 5110 -26174 5170 -25968
rect 5110 -26240 5170 -26234
rect 6132 -26174 6192 -25968
rect 6132 -26240 6192 -26234
rect 6640 -26430 6700 -25204
rect 7154 -25294 7214 -25094
rect 8168 -25284 8228 -25094
rect 8678 -25144 8738 -24686
rect 9694 -24686 9706 -24660
rect 9740 -24592 9746 -24110
rect 10712 -24110 10772 -23882
rect 11006 -24026 11218 -24020
rect 11278 -24026 11494 -24020
rect 11006 -24060 11018 -24026
rect 11482 -24060 11494 -24026
rect 11006 -24066 11494 -24060
rect 12024 -24026 12228 -24020
rect 12288 -24026 12512 -24020
rect 12024 -24060 12036 -24026
rect 12500 -24060 12512 -24026
rect 12024 -24066 12512 -24060
rect 12742 -24110 12802 -23882
rect 13042 -24026 13242 -24020
rect 13302 -24026 13530 -24020
rect 13042 -24060 13054 -24026
rect 13518 -24060 13530 -24026
rect 13042 -24066 13530 -24060
rect 14060 -24026 14270 -24020
rect 14330 -24026 14548 -24020
rect 14060 -24060 14072 -24026
rect 14536 -24060 14548 -24026
rect 14060 -24066 14548 -24060
rect 14780 -24110 14840 -23882
rect 15078 -24026 15566 -24020
rect 15078 -24060 15090 -24026
rect 15554 -24060 15566 -24026
rect 15078 -24066 15566 -24060
rect 16096 -24026 16584 -24020
rect 16096 -24060 16108 -24026
rect 16572 -24060 16584 -24026
rect 16096 -24066 16584 -24060
rect 10712 -24166 10724 -24110
rect 10718 -24592 10724 -24166
rect 9740 -24686 9754 -24660
rect 9200 -25034 9260 -24770
rect 9694 -24928 9754 -24686
rect 10716 -24686 10724 -24662
rect 10758 -24166 10772 -24110
rect 11730 -24146 11742 -24110
rect 10758 -24592 10764 -24166
rect 11736 -24592 11742 -24146
rect 10758 -24686 10776 -24662
rect 10212 -24736 10272 -24734
rect 9842 -24882 9848 -24822
rect 9908 -24882 9914 -24822
rect 9688 -24988 9694 -24928
rect 9754 -24988 9760 -24928
rect 9194 -25094 9200 -25034
rect 9260 -25094 9266 -25034
rect 9848 -25066 9908 -24882
rect 10212 -25034 10272 -24770
rect 8672 -25204 8678 -25144
rect 8738 -25204 8744 -25144
rect 7144 -26168 7204 -25964
rect 7654 -26066 7714 -25876
rect 7648 -26126 7654 -26066
rect 7714 -26126 7720 -26066
rect 8170 -26168 8230 -25964
rect 7144 -26174 7206 -26168
rect 7144 -26180 7146 -26174
rect 8170 -26174 8232 -26168
rect 8170 -26180 8172 -26174
rect 7146 -26240 7206 -26234
rect 8172 -26240 8232 -26234
rect 8678 -26430 8738 -25204
rect 9200 -25290 9260 -25094
rect 9692 -25126 9908 -25066
rect 10206 -25094 10212 -25034
rect 10272 -25094 10278 -25034
rect 9692 -25368 9752 -25126
rect 10212 -25288 10272 -25094
rect 10716 -25144 10776 -24686
rect 11726 -24686 11742 -24634
rect 11776 -24146 11790 -24110
rect 11776 -24592 11782 -24146
rect 12742 -24160 12760 -24110
rect 12754 -24592 12760 -24160
rect 11776 -24686 11786 -24634
rect 11220 -25034 11280 -24770
rect 11726 -24822 11786 -24686
rect 12752 -24686 12760 -24656
rect 12794 -24160 12802 -24110
rect 13766 -24142 13778 -24110
rect 12794 -24592 12800 -24160
rect 13772 -24592 13778 -24142
rect 12794 -24686 12812 -24656
rect 11720 -24882 11726 -24822
rect 11786 -24882 11792 -24822
rect 11724 -24988 11730 -24928
rect 11790 -24988 11796 -24928
rect 11214 -25094 11220 -25034
rect 11280 -25094 11286 -25034
rect 10710 -25204 10716 -25144
rect 10776 -25204 10782 -25144
rect 9184 -26174 9244 -25968
rect 9184 -26240 9244 -26234
rect 10220 -26174 10280 -25972
rect 10220 -26240 10280 -26234
rect 10716 -26430 10776 -25204
rect 11220 -25290 11280 -25094
rect 11730 -25368 11790 -24988
rect 12238 -25034 12298 -24770
rect 12232 -25094 12238 -25034
rect 12298 -25094 12304 -25034
rect 12238 -25288 12298 -25094
rect 12752 -25144 12812 -24686
rect 13764 -24686 13778 -24646
rect 13812 -24142 13826 -24110
rect 13812 -24592 13818 -24142
rect 14780 -24154 14796 -24110
rect 14790 -24592 14796 -24154
rect 13812 -24686 13824 -24646
rect 13264 -25034 13324 -24770
rect 13764 -24822 13824 -24686
rect 14788 -24686 14796 -24662
rect 14830 -24154 14840 -24110
rect 15808 -24110 15854 -24098
rect 14830 -24592 14836 -24154
rect 15808 -24592 15814 -24110
rect 14830 -24686 14848 -24662
rect 13758 -24882 13764 -24822
rect 13824 -24882 13830 -24822
rect 13760 -24988 13766 -24928
rect 13826 -24988 13832 -24928
rect 13258 -25094 13264 -25034
rect 13324 -25094 13330 -25034
rect 12746 -25204 12752 -25144
rect 12812 -25204 12818 -25144
rect 11226 -26174 11286 -25972
rect 12240 -26174 12300 -25972
rect 12234 -26234 12240 -26174
rect 12300 -26234 12306 -26174
rect 11226 -26240 11286 -26234
rect 12752 -26430 12812 -25204
rect 13264 -25288 13324 -25094
rect 13766 -25378 13826 -24988
rect 14266 -25034 14326 -24770
rect 14260 -25094 14266 -25034
rect 14326 -25094 14332 -25034
rect 14266 -25290 14326 -25094
rect 14788 -25144 14848 -24686
rect 15800 -24686 15814 -24640
rect 15848 -24592 15854 -24110
rect 16816 -24110 16876 -23882
rect 16962 -23926 17022 -23662
rect 16956 -23986 16962 -23926
rect 17022 -23986 17028 -23926
rect 17326 -24020 17386 -23542
rect 17838 -23822 17898 -23452
rect 18856 -23452 18868 -23408
rect 18902 -23408 18908 -22876
rect 19870 -22876 19930 -22738
rect 20396 -22786 20456 -22736
rect 21410 -22786 21470 -22608
rect 21904 -22736 21910 -22676
rect 21970 -22736 21976 -22676
rect 20168 -22792 20656 -22786
rect 20168 -22826 20180 -22792
rect 20644 -22826 20656 -22792
rect 20168 -22832 20656 -22826
rect 21186 -22792 21674 -22786
rect 21186 -22826 21198 -22792
rect 21662 -22826 21674 -22792
rect 21186 -22832 21674 -22826
rect 19870 -22922 19886 -22876
rect 19880 -23404 19886 -22922
rect 18902 -23452 18916 -23408
rect 18132 -23502 18620 -23496
rect 18132 -23536 18144 -23502
rect 18608 -23536 18620 -23502
rect 18132 -23542 18620 -23536
rect 17832 -23882 17838 -23822
rect 17898 -23882 17904 -23822
rect 18346 -24020 18406 -23542
rect 18856 -23594 18916 -23452
rect 19872 -23452 19886 -23404
rect 19920 -22922 19930 -22876
rect 20898 -22876 20944 -22864
rect 21910 -22876 21970 -22736
rect 22204 -22792 22410 -22786
rect 22470 -22792 22692 -22786
rect 22204 -22826 22216 -22792
rect 22680 -22826 22692 -22792
rect 22204 -22832 22692 -22826
rect 19920 -23404 19926 -22922
rect 19920 -23452 19932 -23404
rect 20898 -23408 20904 -22876
rect 19150 -23502 19638 -23496
rect 19150 -23536 19162 -23502
rect 19626 -23536 19638 -23502
rect 19150 -23542 19638 -23536
rect 18850 -23654 18856 -23594
rect 18916 -23654 18922 -23594
rect 18852 -23882 18858 -23822
rect 18918 -23882 18924 -23822
rect 17114 -24026 17602 -24020
rect 17114 -24060 17126 -24026
rect 17590 -24060 17602 -24026
rect 17114 -24066 17602 -24060
rect 18132 -24026 18620 -24020
rect 18132 -24060 18144 -24026
rect 18608 -24060 18620 -24026
rect 18132 -24066 18620 -24060
rect 16816 -24154 16832 -24110
rect 16826 -24592 16832 -24154
rect 15848 -24686 15860 -24640
rect 15286 -25034 15346 -24770
rect 15628 -24882 15634 -24822
rect 15694 -24882 15700 -24822
rect 15280 -25094 15286 -25034
rect 15346 -25094 15352 -25034
rect 15634 -25074 15694 -24882
rect 15800 -24928 15860 -24686
rect 16820 -24686 16832 -24660
rect 16866 -24154 16876 -24110
rect 17844 -24110 17890 -24098
rect 16866 -24592 16872 -24154
rect 17844 -24592 17850 -24110
rect 16866 -24686 16880 -24660
rect 15794 -24988 15800 -24928
rect 15860 -24988 15866 -24928
rect 16306 -25034 16366 -24770
rect 14782 -25204 14788 -25144
rect 14848 -25204 14854 -25144
rect 13256 -26174 13316 -25968
rect 14266 -26168 14326 -25972
rect 13256 -26240 13316 -26234
rect 14264 -26174 14326 -26168
rect 14324 -26180 14326 -26174
rect 14264 -26240 14324 -26234
rect 14788 -26430 14848 -25204
rect 15286 -25288 15346 -25094
rect 15634 -25134 15860 -25074
rect 16300 -25094 16306 -25034
rect 16366 -25094 16372 -25034
rect 15800 -25378 15860 -25134
rect 16306 -25288 16366 -25094
rect 16820 -25144 16880 -24686
rect 17840 -24686 17850 -24646
rect 17884 -24592 17890 -24110
rect 18858 -24110 18918 -23882
rect 19360 -24020 19420 -23542
rect 19872 -23822 19932 -23452
rect 20888 -23452 20904 -23408
rect 20938 -23408 20944 -22876
rect 21908 -22910 21922 -22876
rect 21910 -22920 21922 -22910
rect 20938 -23452 20948 -23408
rect 20168 -23502 20656 -23496
rect 20168 -23536 20180 -23502
rect 20644 -23536 20656 -23502
rect 20168 -23542 20656 -23536
rect 19866 -23882 19872 -23822
rect 19932 -23882 19938 -23822
rect 19866 -23986 19872 -23926
rect 19932 -23986 19938 -23926
rect 19150 -24026 19420 -24020
rect 19428 -24026 19638 -24020
rect 19150 -24060 19162 -24026
rect 19626 -24060 19638 -24026
rect 19150 -24066 19638 -24060
rect 19368 -24070 19428 -24066
rect 18858 -24176 18868 -24110
rect 18862 -24592 18868 -24176
rect 17884 -24686 17900 -24646
rect 17332 -25034 17392 -24770
rect 17840 -24928 17900 -24686
rect 18852 -24686 18868 -24640
rect 18902 -24176 18918 -24110
rect 19872 -24110 19932 -23986
rect 20396 -24020 20456 -23542
rect 20888 -23594 20948 -23452
rect 21916 -23452 21922 -22920
rect 21956 -22920 21970 -22876
rect 22922 -22876 22982 -22608
rect 21956 -23452 21962 -22920
rect 22922 -22930 22940 -22876
rect 21916 -23464 21962 -23452
rect 22934 -23452 22940 -22930
rect 22974 -22914 22986 -22876
rect 22974 -22930 22982 -22914
rect 22974 -23452 22980 -22930
rect 22934 -23464 22980 -23452
rect 21186 -23502 21674 -23496
rect 21186 -23536 21198 -23502
rect 21662 -23536 21674 -23502
rect 21186 -23542 21674 -23536
rect 22204 -23502 22692 -23496
rect 22204 -23536 22216 -23502
rect 22680 -23536 22692 -23502
rect 22204 -23542 22692 -23536
rect 20882 -23654 20888 -23594
rect 20948 -23654 20954 -23594
rect 21408 -23704 21468 -23542
rect 22416 -23704 22476 -23542
rect 23034 -23594 23094 -17804
rect 23156 -18718 23162 -18658
rect 23222 -18718 23228 -18658
rect 23162 -20216 23222 -18718
rect 23278 -18982 23338 -17690
rect 23394 -18940 23400 -18880
rect 23460 -18940 23466 -18880
rect 23272 -19042 23278 -18982
rect 23338 -19042 23344 -18982
rect 23156 -20276 23162 -20216
rect 23222 -20276 23228 -20216
rect 23152 -21178 23158 -21118
rect 23218 -21178 23224 -21118
rect 23158 -22442 23218 -21178
rect 23278 -22344 23338 -19042
rect 23272 -22404 23278 -22344
rect 23338 -22404 23344 -22344
rect 23152 -22502 23158 -22442
rect 23218 -22502 23224 -22442
rect 23028 -23654 23034 -23594
rect 23094 -23654 23100 -23594
rect 21402 -23764 21408 -23704
rect 21468 -23764 21474 -23704
rect 22410 -23764 22416 -23704
rect 22476 -23764 22482 -23704
rect 23278 -23820 23338 -22404
rect 23400 -22676 23460 -18940
rect 23528 -20108 23588 -17586
rect 23526 -20114 23588 -20108
rect 23586 -20174 23588 -20114
rect 23526 -20180 23588 -20174
rect 23528 -22548 23588 -20180
rect 23522 -22608 23528 -22548
rect 23588 -22608 23594 -22548
rect 23394 -22736 23400 -22676
rect 23460 -22736 23466 -22676
rect 23650 -23704 23710 -12776
rect 23756 -16586 23762 -16526
rect 23822 -16586 23828 -16526
rect 23644 -23764 23650 -23704
rect 23710 -23764 23716 -23704
rect 20888 -23882 20894 -23822
rect 20954 -23882 20960 -23822
rect 21910 -23880 23338 -23820
rect 20168 -24026 20656 -24020
rect 20168 -24060 20180 -24026
rect 20644 -24060 20656 -24026
rect 20168 -24066 20656 -24060
rect 19872 -24156 19886 -24110
rect 18902 -24592 18908 -24176
rect 19880 -24592 19886 -24156
rect 18902 -24686 18912 -24640
rect 19920 -24156 19932 -24110
rect 20894 -24110 20954 -23882
rect 21186 -24026 21408 -24020
rect 21468 -24026 21674 -24020
rect 21186 -24060 21198 -24026
rect 21662 -24060 21674 -24026
rect 21186 -24066 21674 -24060
rect 19920 -24592 19926 -24156
rect 20894 -24170 20904 -24110
rect 20898 -24592 20904 -24170
rect 20892 -24686 20904 -24662
rect 20938 -24170 20954 -24110
rect 21910 -24110 21970 -23880
rect 22408 -24020 22468 -23880
rect 22204 -24026 22692 -24020
rect 22204 -24060 22216 -24026
rect 22680 -24060 22692 -24026
rect 22204 -24066 22692 -24060
rect 20938 -24592 20944 -24170
rect 20938 -24686 20952 -24662
rect 18350 -24736 18410 -24734
rect 17834 -24988 17840 -24928
rect 17900 -24988 17906 -24928
rect 18350 -25034 18410 -24770
rect 17326 -25094 17332 -25034
rect 17392 -25094 17398 -25034
rect 18344 -25094 18350 -25034
rect 18410 -25094 18416 -25034
rect 16814 -25204 16820 -25144
rect 16880 -25204 16886 -25144
rect 15282 -26168 15342 -25972
rect 15280 -26174 15342 -26168
rect 15340 -26180 15342 -26174
rect 16304 -26174 16364 -25960
rect 15280 -26240 15340 -26234
rect 16304 -26240 16364 -26234
rect 16820 -26430 16880 -25204
rect 17332 -25294 17392 -25094
rect 18350 -25294 18410 -25094
rect 18852 -25144 18912 -24686
rect 19364 -25034 19424 -24770
rect 19864 -24988 19870 -24928
rect 19930 -24988 19936 -24928
rect 19358 -25094 19364 -25034
rect 19424 -25094 19430 -25034
rect 18846 -25204 18852 -25144
rect 18912 -25204 18918 -25144
rect 17326 -26174 17386 -25964
rect 17834 -26066 17894 -25866
rect 17828 -26126 17834 -26066
rect 17894 -26126 17900 -26066
rect 18346 -26168 18406 -25972
rect 18346 -26174 18408 -26168
rect 18346 -26180 18348 -26174
rect 17326 -26240 17386 -26234
rect 18348 -26240 18408 -26234
rect 18852 -26430 18912 -25204
rect 19364 -25284 19424 -25094
rect 19870 -25386 19930 -24988
rect 20378 -25034 20438 -24770
rect 20372 -25094 20378 -25034
rect 20438 -25094 20444 -25034
rect 20378 -25284 20438 -25094
rect 20892 -25144 20952 -24686
rect 21910 -24686 21922 -24110
rect 21956 -24686 21970 -24110
rect 22924 -24110 22984 -23880
rect 23048 -23986 23054 -23926
rect 23114 -23986 23120 -23926
rect 22924 -24164 22940 -24110
rect 22934 -24592 22940 -24164
rect 22974 -24164 22984 -24110
rect 22974 -24592 22980 -24164
rect 21400 -24736 21460 -24734
rect 21400 -25034 21460 -24770
rect 21910 -24822 21970 -24686
rect 21904 -24882 21910 -24822
rect 21970 -24882 21976 -24822
rect 21904 -24988 21910 -24928
rect 21970 -24988 21976 -24928
rect 21394 -25094 21400 -25034
rect 21460 -25094 21466 -25034
rect 20886 -25204 20892 -25144
rect 20952 -25204 20958 -25144
rect 19368 -26168 19428 -25960
rect 20382 -26168 20442 -25968
rect 19366 -26174 19428 -26168
rect 19426 -26180 19428 -26174
rect 20380 -26174 20442 -26168
rect 19366 -26240 19426 -26234
rect 20440 -26180 20442 -26174
rect 20380 -26240 20440 -26234
rect 20892 -26430 20952 -25204
rect 21400 -25284 21460 -25094
rect 21910 -25144 21970 -24988
rect 21910 -25204 22988 -25144
rect 21910 -25350 21970 -25204
rect 22426 -25294 22486 -25204
rect 22928 -25360 22988 -25204
rect 21402 -26168 21462 -25960
rect 23054 -26066 23114 -23986
rect 23762 -24928 23822 -16586
rect 23756 -24988 23762 -24928
rect 23822 -24988 23828 -24928
rect 23048 -26126 23054 -26066
rect 23114 -26126 23120 -26066
rect 21402 -26174 21464 -26168
rect 21402 -26180 21404 -26174
rect 21404 -26240 21464 -26234
rect 24816 -26330 24822 -12070
rect 24922 -26330 24928 -12070
rect -8118 -26476 -7968 -26430
rect -7922 -26476 -4748 -26430
rect -4688 -26476 1704 -26430
rect 1764 -26476 23806 -26430
rect 23866 -26476 23968 -26430
rect -8118 -26630 -8072 -26476
rect 23928 -26630 23968 -26476
rect -8118 -26676 23968 -26630
rect -11616 -27116 -11606 -26816
rect 24206 -27116 24216 -26816
rect 24816 -27116 24928 -26330
rect -12328 -27122 24928 -27116
rect -12328 -27222 -12222 -27122
rect 24822 -27222 24928 -27122
rect -12328 -27228 24928 -27222
<< via1 >>
rect 484 3916 1084 4216
rect 24116 3916 24716 4216
rect 4061 3620 20846 3834
rect 7986 1858 8046 1918
rect 9068 1858 9128 1918
rect 10026 1858 10086 1918
rect 8512 1612 8572 1672
rect 10548 1612 10608 1672
rect 13090 1858 13150 1918
rect 14108 1858 14168 1918
rect 12586 1614 12646 1674
rect 15132 1858 15192 1918
rect 16144 1858 16204 1918
rect 14616 1614 14676 1674
rect 16658 1616 16718 1676
rect 17668 1616 17728 1676
rect 19202 1858 19262 1918
rect 20214 1858 20274 1918
rect 18690 1616 18750 1676
rect 21232 1858 21292 1918
rect 20726 1616 20786 1676
rect 6330 680 6390 740
rect 7494 680 7554 740
rect 6200 476 6260 536
rect 4192 -1708 4252 -1648
rect 3676 -5966 3736 -5906
rect 3784 -6078 3844 -6018
rect 2014 -7000 2074 -6940
rect 3174 -7110 3234 -7050
rect 1888 -8088 1948 -8028
rect 3690 -8034 3750 -7974
rect 3796 -8134 3856 -8074
rect 7494 476 7554 536
rect 9530 576 9590 636
rect 11566 576 11626 636
rect 13604 680 13664 740
rect 13600 476 13660 536
rect 15638 680 15698 740
rect 15636 476 15696 536
rect 16138 476 16198 536
rect 17672 576 17732 636
rect 17158 476 17218 536
rect 18184 476 18244 536
rect 19706 576 19766 636
rect 18690 472 18750 532
rect 19204 472 19264 532
rect 19708 472 19768 532
rect 20214 472 20274 532
rect 20734 472 20794 532
rect 21746 680 21806 740
rect 22996 680 23056 740
rect 7980 -674 8040 -614
rect 10036 -458 10096 -398
rect 10546 -458 10606 -398
rect 9528 -560 9592 -496
rect 9018 -674 9078 -614
rect 10030 -674 10090 -614
rect 11404 -560 11468 -496
rect 12580 -458 12640 -398
rect 11040 -666 11100 -606
rect 12064 -666 12124 -606
rect 13092 -666 13152 -606
rect 14618 -460 14678 -400
rect 15638 -558 15698 -498
rect 16654 -460 16714 -400
rect 17154 -460 17214 -400
rect 17668 -460 17728 -400
rect 18192 -460 18252 -400
rect 18690 -460 18750 -400
rect 19192 -460 19252 -400
rect 19706 -462 19766 -402
rect 20214 -462 20274 -402
rect 20724 -462 20784 -402
rect 19196 -674 19256 -614
rect 20208 -674 20268 -614
rect 21746 -558 21806 -498
rect 21210 -674 21270 -614
rect 6330 -1994 6390 -1934
rect 6686 -4402 6746 -4342
rect 6560 -5012 6620 -4952
rect 4698 -5966 4758 -5906
rect 4568 -6078 4628 -6018
rect 5208 -7000 5268 -6940
rect 6360 -7110 6420 -7050
rect 4700 -8034 4760 -7974
rect 6552 -7238 6612 -7178
rect 4582 -8134 4642 -8074
rect 1402 -9144 1462 -9084
rect 1542 -9320 1602 -9260
rect 2442 -9494 2502 -9434
rect 6802 -5012 6862 -4952
rect 7488 -1848 7552 -1784
rect 7312 -1994 7372 -1934
rect 8510 -1596 8570 -1536
rect 9526 -1710 9590 -1646
rect 10546 -1596 10606 -1536
rect 11068 -1596 11128 -1536
rect 11566 -1596 11626 -1536
rect 12040 -1600 12100 -1540
rect 7428 -2100 7488 -2040
rect 7990 -2100 8050 -2040
rect 9032 -2100 9092 -2040
rect 10032 -2100 10092 -2040
rect 12580 -1538 12640 -1536
rect 12548 -1596 12640 -1538
rect 13040 -1596 13100 -1536
rect 12548 -1598 12608 -1596
rect 13598 -1852 13662 -1788
rect 14084 -1594 14144 -1534
rect 13194 -2100 13254 -2040
rect 14616 -1596 14676 -1536
rect 16128 -1594 16188 -1534
rect 15634 -1994 15698 -1930
rect 14204 -2100 14264 -2040
rect 15146 -2100 15206 -2040
rect 16654 -1540 16714 -1538
rect 16622 -1598 16714 -1540
rect 16622 -1600 16682 -1598
rect 17150 -1604 17210 -1544
rect 17638 -1542 17698 -1540
rect 17638 -1600 17732 -1542
rect 17672 -1602 17732 -1600
rect 18150 -1604 18210 -1544
rect 18690 -1600 18750 -1540
rect 20724 -1600 20784 -1540
rect 19706 -1710 19770 -1646
rect 22992 -1848 23056 -1784
rect 21740 -1994 21800 -1934
rect 7542 -2302 7602 -2242
rect 8686 -3238 8746 -3178
rect 9190 -3346 9250 -3286
rect 8682 -4270 8742 -4210
rect 9188 -4404 9248 -4344
rect 10720 -2302 10780 -2242
rect 10720 -3238 10780 -3178
rect 10212 -3346 10272 -3286
rect 11230 -3346 11290 -3286
rect 10202 -4408 10262 -4348
rect 11234 -4400 11294 -4340
rect 12762 -3238 12822 -3178
rect 12254 -3346 12314 -3286
rect 13268 -3346 13328 -3286
rect 12762 -4270 12822 -4210
rect 12232 -4400 12292 -4340
rect 13276 -4400 13336 -4340
rect 14788 -2302 14848 -2242
rect 14788 -3238 14848 -3178
rect 14286 -3346 14346 -3286
rect 15296 -3346 15356 -3286
rect 14280 -4404 14340 -4344
rect 15296 -4404 15356 -4344
rect 14080 -4612 14140 -4552
rect 7312 -4930 7372 -4870
rect 8478 -4930 8538 -4870
rect 7044 -5976 7104 -5916
rect 6802 -7134 6862 -7074
rect 6798 -7348 6858 -7288
rect 6686 -8390 6746 -8330
rect 1282 -9644 1342 -9584
rect 7180 -6074 7240 -6014
rect 7044 -9648 7104 -9588
rect 10514 -4930 10574 -4870
rect 11022 -4934 11086 -4870
rect 9496 -5878 9556 -5818
rect 11532 -5878 11592 -5818
rect 11874 -5876 11934 -5816
rect 18864 -2302 18924 -2242
rect 16830 -3238 16890 -3178
rect 16318 -3346 16378 -3286
rect 17332 -3346 17392 -3286
rect 16830 -4270 16890 -4210
rect 16300 -4404 16360 -4344
rect 17332 -4400 17392 -4340
rect 15816 -4612 15876 -4552
rect 15096 -4812 15160 -4748
rect 18866 -3238 18926 -3178
rect 18364 -3346 18424 -3286
rect 19374 -3346 19434 -3286
rect 18348 -4404 18408 -4344
rect 19376 -4404 19436 -4344
rect 22060 -2302 22120 -2242
rect 20902 -3238 20962 -3178
rect 20396 -3346 20456 -3286
rect 20898 -4270 20958 -4210
rect 20396 -4404 20456 -4344
rect 22854 -4402 22914 -4342
rect 21714 -4628 21774 -4568
rect 19160 -4812 19224 -4748
rect 20184 -4812 20248 -4748
rect 21196 -4812 21260 -4748
rect 15098 -4934 15162 -4870
rect 9496 -6074 9556 -6014
rect 10516 -6072 10576 -6012
rect 8482 -6184 8542 -6124
rect 10516 -6184 10576 -6124
rect 14588 -5876 14648 -5816
rect 18660 -4930 18720 -4870
rect 20694 -4930 20754 -4870
rect 15606 -6072 15666 -6012
rect 13572 -6186 13632 -6126
rect 15606 -6186 15666 -6126
rect 18662 -6186 18722 -6126
rect 19676 -5878 19736 -5818
rect 20696 -6186 20756 -6126
rect 21712 -5878 21772 -5818
rect 7464 -7348 7524 -7288
rect 9498 -7238 9558 -7178
rect 9498 -7442 9558 -7382
rect 11534 -7238 11594 -7178
rect 11532 -7340 11592 -7280
rect 11532 -7442 11592 -7382
rect 13568 -7134 13628 -7074
rect 14588 -7134 14648 -7074
rect 14588 -7440 14648 -7380
rect 15606 -7440 15666 -7380
rect 16624 -7134 16684 -7074
rect 16622 -7440 16682 -7380
rect 18658 -7238 18718 -7178
rect 19526 -7120 19586 -7060
rect 19674 -7230 19734 -7170
rect 19526 -7440 19586 -7380
rect 19678 -7438 19738 -7378
rect 20694 -7340 20754 -7280
rect 23290 -4270 23350 -4210
rect 22996 -4630 23056 -4570
rect 23138 -4930 23198 -4870
rect 22978 -6072 23038 -6012
rect 21714 -7230 21774 -7170
rect 22854 -7230 22914 -7170
rect 21712 -7438 21772 -7378
rect 8480 -8390 8540 -8330
rect 7312 -8598 7372 -8538
rect 9494 -8700 9554 -8640
rect 10516 -8390 10576 -8330
rect 10516 -8498 10576 -8438
rect 11534 -8382 11594 -8322
rect 13336 -8382 13396 -8322
rect 11528 -8700 11588 -8640
rect 11732 -8712 11792 -8652
rect 13570 -8388 13630 -8328
rect 15606 -8388 15666 -8328
rect 15604 -8498 15664 -8438
rect 15094 -8712 15154 -8652
rect 16110 -8712 16170 -8652
rect 18660 -8386 18720 -8326
rect 19170 -8712 19230 -8652
rect 19682 -8700 19742 -8640
rect 20696 -8386 20756 -8326
rect 22978 -7438 23038 -7378
rect 22854 -8498 22914 -8438
rect 21716 -8700 21776 -8640
rect 8476 -9648 8536 -9588
rect 10512 -9648 10572 -9588
rect 7180 -9778 7240 -9718
rect 2336 -9906 2396 -9846
rect 2216 -10024 2276 -9964
rect 18664 -9648 18724 -9588
rect 20700 -9648 20760 -9588
rect 11534 -9918 11594 -9858
rect 23290 -6186 23350 -6126
rect 23138 -9918 23198 -9858
rect 1770 -10142 1830 -10082
rect -13630 -10670 -2866 -10378
rect 1888 -11418 1948 -11358
rect 2216 -11408 2276 -11348
rect 1282 -11554 1342 -11494
rect 1402 -11552 1462 -11492
rect 1542 -11534 1602 -11474
rect 1770 -11518 1830 -11458
rect 1150 -11682 1210 -11622
rect -1562 -12280 -1502 -12220
rect -36 -12414 24 -12354
rect 1150 -18882 1210 -18822
rect -3398 -19808 -3338 -19748
rect -9508 -19954 -9448 -19894
rect -5428 -19954 -5368 -19894
rect -10662 -20082 -10602 -20022
rect -7984 -20082 -7924 -20022
rect -6952 -20082 -6892 -20022
rect -3892 -20082 -3832 -20022
rect -9004 -21044 -8944 -20984
rect -9504 -21148 -9444 -21088
rect -10662 -22314 -10602 -22254
rect -7980 -21044 -7920 -20984
rect -8486 -21252 -8426 -21192
rect -9012 -22314 -8952 -22254
rect -6948 -21044 -6888 -20984
rect -7468 -21148 -7408 -21088
rect -5948 -21044 -5888 -20984
rect -4928 -21044 -4868 -20984
rect -5432 -21148 -5372 -21088
rect -6450 -21252 -6390 -21192
rect -7474 -22194 -7414 -22134
rect -8486 -23258 -8426 -23198
rect -9500 -23366 -9440 -23306
rect -9006 -23478 -8946 -23418
rect -7464 -23366 -7404 -23306
rect -7982 -23478 -7922 -23418
rect -5942 -22314 -5882 -22254
rect -3908 -21044 -3848 -20984
rect -4418 -21252 -4358 -21192
rect -4934 -22314 -4874 -22254
rect -6450 -23258 -6390 -23198
rect -6950 -23478 -6890 -23418
rect -1368 -19954 -1308 -19894
rect 816 -19954 876 -19894
rect -2896 -20082 -2836 -20022
rect -2898 -21044 -2838 -20984
rect -3398 -21148 -3338 -21088
rect -1884 -21044 -1824 -20984
rect -866 -21044 -806 -20984
rect -1362 -21148 -1302 -21088
rect -2384 -21252 -2324 -21192
rect -3398 -22194 -3338 -22134
rect -4418 -23258 -4358 -23198
rect -5428 -23366 -5368 -23306
rect -5950 -23478 -5890 -23418
rect -4930 -23478 -4870 -23418
rect -3394 -23366 -3334 -23306
rect -3910 -23478 -3850 -23418
rect -2900 -23478 -2840 -23418
rect -1872 -22314 -1812 -22254
rect -340 -21252 -280 -21192
rect 936 -21044 996 -20984
rect 816 -22194 876 -22134
rect -846 -22314 -786 -22254
rect -2384 -23258 -2324 -23198
rect -340 -23258 -280 -23198
rect -1358 -23366 -1298 -23306
rect -1886 -23478 -1826 -23418
rect -868 -23478 -808 -23418
rect -10662 -24440 -10602 -24380
rect -7992 -24440 -7932 -24380
rect -6960 -24440 -6900 -24380
rect -3900 -24440 -3840 -24380
rect -2904 -24440 -2844 -24380
rect 936 -23478 996 -23418
rect -9506 -24570 -9446 -24510
rect -5426 -24570 -5366 -24510
rect -1366 -24570 -1306 -24510
rect 816 -24570 876 -24510
rect -8028 -25936 -7968 -25876
rect -5990 -25936 -5930 -25876
rect -3954 -25936 -3894 -25876
rect -7010 -26048 -6950 -25988
rect -1918 -25936 -1858 -25876
rect -2936 -26048 -2876 -25988
rect 1282 -19954 1342 -19894
rect 1402 -20082 1462 -20022
rect 1660 -11672 1720 -11612
rect 1770 -12414 1830 -12354
rect 2336 -11416 2396 -11356
rect 2216 -12280 2276 -12220
rect 2012 -13638 2072 -13578
rect 1886 -15340 1946 -15280
rect 1660 -17800 1720 -17740
rect 1542 -21044 1602 -20984
rect 2224 -13974 2284 -13914
rect 2120 -15234 2180 -15174
rect 2012 -16334 2072 -16274
rect 2442 -11552 2502 -11492
rect 13254 -11902 13314 -11842
rect 18358 -11902 18418 -11842
rect 22418 -11908 22478 -11848
rect 3586 -13638 3646 -13578
rect 4600 -13854 4660 -13794
rect 6640 -13854 6700 -13794
rect 8680 -13854 8740 -13794
rect 10710 -13854 10770 -13794
rect 12750 -13854 12810 -13794
rect 14782 -13854 14842 -13794
rect 16822 -13854 16882 -13794
rect 18858 -13854 18918 -13794
rect 20892 -13854 20952 -13794
rect 2568 -13974 2628 -13914
rect 4092 -13980 4152 -13920
rect 2442 -14096 2502 -14036
rect 5106 -13980 5166 -13920
rect 6128 -13980 6188 -13920
rect 7142 -13980 7202 -13920
rect 8168 -13980 8228 -13920
rect 7656 -14096 7716 -14036
rect 9180 -13980 9240 -13920
rect 10216 -13980 10276 -13920
rect 11222 -13980 11282 -13920
rect 12236 -13980 12296 -13920
rect 13252 -13980 13312 -13920
rect 14260 -13980 14320 -13920
rect 15276 -13980 15336 -13920
rect 16300 -13980 16360 -13920
rect 17322 -13980 17382 -13920
rect 18344 -13980 18404 -13920
rect 17844 -14096 17904 -14036
rect 4604 -15018 4664 -14958
rect 4096 -15128 4156 -15068
rect 3586 -15234 3646 -15174
rect 2572 -15340 2632 -15280
rect 3070 -15340 3130 -15280
rect 3582 -15340 3642 -15280
rect 5118 -15128 5178 -15068
rect 6644 -15018 6704 -14958
rect 6132 -15128 6192 -15068
rect 5626 -15234 5686 -15174
rect 8676 -15018 8736 -14958
rect 7146 -15128 7206 -15068
rect 8164 -15128 8224 -15068
rect 7656 -15234 7716 -15174
rect 2442 -16230 2502 -16170
rect 2566 -16334 2626 -16274
rect 4086 -16334 4146 -16274
rect 4598 -16334 4658 -16274
rect 2336 -16456 2396 -16396
rect 2224 -16570 2284 -16510
rect 3072 -16570 3132 -16510
rect 4604 -16568 4664 -16508
rect 9190 -15128 9250 -15068
rect 10708 -15018 10768 -14958
rect 9696 -15234 9756 -15174
rect 10210 -15128 10270 -15068
rect 9862 -15340 9922 -15280
rect 5620 -16230 5680 -16170
rect 5622 -16334 5682 -16274
rect 11230 -15128 11290 -15068
rect 12744 -15018 12804 -14958
rect 12232 -15128 12292 -15068
rect 11730 -15234 11790 -15174
rect 11730 -15340 11790 -15280
rect 13258 -15128 13318 -15068
rect 19362 -13980 19422 -13920
rect 20376 -13980 20436 -13920
rect 21400 -13980 21460 -13920
rect 21916 -14096 21976 -14036
rect 23048 -14096 23108 -14036
rect 14780 -15018 14840 -14958
rect 14276 -15128 14336 -15068
rect 13766 -15234 13826 -15174
rect 13768 -15340 13828 -15280
rect 15284 -15128 15344 -15068
rect 16818 -15018 16878 -14958
rect 16296 -15128 16356 -15068
rect 15802 -15234 15862 -15174
rect 15648 -15340 15708 -15280
rect 18856 -15018 18916 -14958
rect 17328 -15128 17388 -15068
rect 18342 -15128 18402 -15068
rect 17842 -15234 17902 -15174
rect 6634 -16334 6694 -16274
rect 6640 -16568 6700 -16508
rect 7654 -16334 7714 -16274
rect 2448 -17498 2508 -17438
rect 3586 -17498 3646 -17438
rect 2336 -17698 2396 -17638
rect 2230 -17800 2290 -17740
rect 2120 -21252 2180 -21192
rect 2336 -18934 2396 -18874
rect 1888 -21402 1948 -21342
rect 2230 -21290 2290 -21230
rect 3584 -17698 3644 -17638
rect 4602 -17578 4662 -17518
rect 8676 -16230 8736 -16170
rect 14782 -16230 14842 -16170
rect 10712 -16334 10772 -16274
rect 12750 -16334 12810 -16274
rect 9696 -16456 9756 -16396
rect 11730 -16456 11790 -16396
rect 13760 -16456 13820 -16396
rect 5620 -17474 5680 -17414
rect 5116 -17692 5176 -17632
rect 6642 -17578 6702 -17518
rect 6120 -17692 6180 -17632
rect 3584 -18730 3644 -18670
rect 4090 -18832 4150 -18772
rect 7656 -17474 7716 -17414
rect 7132 -17692 7192 -17632
rect 8674 -17578 8734 -17518
rect 8152 -17692 8212 -17632
rect 8674 -17690 8734 -17630
rect 10708 -17578 10768 -17518
rect 9692 -17800 9752 -17740
rect 5622 -18730 5682 -18670
rect 5620 -18934 5680 -18874
rect 10710 -17690 10770 -17630
rect 11726 -17800 11786 -17740
rect 15800 -16334 15860 -16274
rect 19360 -15128 19420 -15068
rect 20892 -15018 20952 -14958
rect 20384 -15128 20444 -15068
rect 19872 -15234 19932 -15174
rect 19872 -15338 19932 -15278
rect 16818 -16334 16878 -16274
rect 17838 -16334 17898 -16274
rect 12748 -17578 12808 -17518
rect 12746 -17690 12806 -17630
rect 14782 -17578 14842 -17518
rect 14978 -17582 15038 -17522
rect 13766 -17800 13826 -17740
rect 14782 -17690 14842 -17630
rect 21404 -15128 21464 -15068
rect 21912 -15234 21972 -15174
rect 23048 -15338 23108 -15278
rect 19876 -16230 19936 -16170
rect 18854 -16334 18914 -16274
rect 20890 -16334 20950 -16274
rect 15800 -17474 15860 -17414
rect 14978 -17800 15038 -17740
rect 15272 -17798 15332 -17738
rect 7658 -18730 7718 -18670
rect 4604 -19034 4664 -18974
rect 6128 -18940 6188 -18880
rect 7150 -18940 7210 -18880
rect 6638 -19034 6698 -18974
rect 9690 -18730 9750 -18670
rect 9182 -18832 9242 -18772
rect 8164 -18940 8224 -18880
rect 9182 -18940 9242 -18880
rect 8674 -19034 8734 -18974
rect 4086 -19958 4146 -19898
rect 4996 -19958 5056 -19898
rect 4086 -20174 4146 -20114
rect 2450 -20278 2510 -20218
rect 5998 -19958 6058 -19898
rect 5124 -20174 5184 -20114
rect 7150 -19958 7210 -19898
rect 6638 -20060 6698 -20000
rect 6138 -20174 6198 -20114
rect 4084 -21186 4144 -21126
rect 3586 -21290 3646 -21230
rect 3582 -21500 3642 -21440
rect 5092 -21186 5152 -21126
rect 4602 -21402 4662 -21342
rect 10202 -18940 10262 -18880
rect 16816 -17690 16876 -17630
rect 16300 -17798 16360 -17738
rect 16818 -17804 16878 -17744
rect 17836 -17474 17896 -17414
rect 18854 -17690 18914 -17630
rect 19870 -17582 19930 -17522
rect 20374 -17586 20434 -17526
rect 23034 -16568 23094 -16508
rect 20894 -17690 20954 -17630
rect 18854 -17804 18914 -17744
rect 14272 -18718 14332 -18658
rect 13766 -18846 13826 -18786
rect 15802 -19044 15862 -18984
rect 8160 -19958 8220 -19898
rect 9166 -19958 9226 -19898
rect 10210 -19958 10270 -19898
rect 10710 -19952 10770 -19892
rect 9164 -20174 9224 -20114
rect 10204 -20174 10264 -20114
rect 9688 -20278 9748 -20218
rect 6106 -21186 6166 -21126
rect 7144 -21186 7204 -21126
rect 6640 -21402 6700 -21342
rect 5620 -21500 5680 -21440
rect 11218 -20174 11278 -20114
rect 12746 -19952 12806 -19892
rect 12226 -20174 12286 -20114
rect 13270 -20174 13330 -20114
rect 11730 -20278 11790 -20218
rect 20892 -17804 20952 -17744
rect 17314 -18940 17374 -18880
rect 14782 -19952 14842 -19892
rect 14260 -20174 14320 -20114
rect 15278 -20174 15338 -20114
rect 13768 -20278 13828 -20218
rect 21910 -17474 21970 -17414
rect 22928 -17456 22988 -17396
rect 23162 -16586 23222 -16526
rect 23528 -17586 23588 -17526
rect 23278 -17690 23338 -17630
rect 19366 -18718 19426 -18658
rect 19504 -18714 19564 -18654
rect 23034 -17804 23094 -17744
rect 20386 -18714 20446 -18654
rect 21392 -18714 21452 -18654
rect 18344 -18940 18404 -18880
rect 19504 -18940 19564 -18880
rect 19872 -18940 19932 -18880
rect 19872 -19044 19932 -18984
rect 21910 -18718 21970 -18658
rect 21910 -18846 21970 -18786
rect 20888 -19042 20948 -18982
rect 16820 -19952 16880 -19892
rect 16812 -20060 16872 -20000
rect 16312 -20174 16372 -20114
rect 15802 -20278 15862 -20218
rect 16314 -20282 16374 -20222
rect 17336 -20282 17396 -20222
rect 17836 -20276 17896 -20216
rect 8162 -21186 8222 -21126
rect 8678 -21180 8738 -21120
rect 10714 -21180 10774 -21120
rect 12746 -21180 12806 -21120
rect 14780 -21180 14840 -21120
rect 7660 -21500 7720 -21440
rect 2448 -22522 2508 -22462
rect 3588 -22738 3648 -22678
rect 4602 -22424 4662 -22364
rect 4606 -22618 4666 -22558
rect 5620 -22522 5680 -22462
rect 11730 -21290 11790 -21230
rect 13766 -21290 13826 -21230
rect 10712 -21402 10772 -21342
rect 9696 -21500 9756 -21440
rect 6638 -22424 6698 -22364
rect 7144 -22522 7204 -22462
rect 6642 -22618 6702 -22558
rect 8676 -22424 8736 -22364
rect 8166 -22522 8226 -22462
rect 7656 -22738 7716 -22678
rect 2336 -23654 2396 -23594
rect 2230 -23780 2290 -23720
rect 9188 -22522 9248 -22462
rect 8670 -22618 8730 -22558
rect 18856 -19952 18916 -19892
rect 18852 -20060 18912 -20000
rect 19344 -20174 19404 -20114
rect 20894 -19952 20954 -19892
rect 20890 -20060 20950 -20000
rect 20382 -20174 20442 -20114
rect 19870 -20276 19930 -20216
rect 15802 -21178 15862 -21118
rect 16156 -21178 16216 -21118
rect 15798 -21290 15858 -21230
rect 15308 -21388 15368 -21328
rect 10538 -22404 10598 -22344
rect 10708 -22404 10768 -22344
rect 10192 -22522 10252 -22462
rect 9690 -22738 9750 -22678
rect 5620 -23780 5680 -23720
rect 6140 -23768 6200 -23708
rect 4602 -23882 4662 -23822
rect 6638 -23882 6698 -23822
rect 5620 -23986 5680 -23926
rect 2448 -24884 2508 -24824
rect 2120 -24988 2180 -24928
rect 3584 -24988 3644 -24928
rect 4092 -25094 4152 -25034
rect 1070 -26048 1130 -25988
rect 10538 -22618 10598 -22558
rect 10714 -22612 10774 -22552
rect 16346 -21388 16406 -21328
rect 17322 -21388 17382 -21328
rect 16156 -21496 16216 -21436
rect 21408 -20174 21468 -20114
rect 21912 -20276 21972 -20216
rect 19874 -21178 19934 -21118
rect 18338 -21388 18398 -21328
rect 20364 -21388 20424 -21328
rect 17836 -21500 17896 -21440
rect 19872 -21500 19932 -21440
rect 12750 -22404 12810 -22344
rect 14782 -22404 14842 -22344
rect 16822 -22404 16882 -22344
rect 15800 -22502 15860 -22442
rect 12742 -22612 12802 -22552
rect 7658 -23882 7718 -23822
rect 8674 -23882 8734 -23822
rect 5618 -24884 5678 -24824
rect 5624 -24988 5684 -24928
rect 5112 -25094 5172 -25034
rect 4604 -25204 4664 -25144
rect 2448 -26126 2508 -26066
rect 3584 -26126 3644 -26066
rect 4096 -26234 4156 -26174
rect 6136 -25094 6196 -25034
rect 9694 -23882 9754 -23822
rect 14786 -22612 14846 -22552
rect 16814 -22612 16874 -22552
rect 17840 -22738 17900 -22678
rect 21394 -21388 21454 -21328
rect 21908 -21500 21968 -21440
rect 18852 -22612 18912 -22552
rect 21906 -22502 21966 -22442
rect 20892 -22612 20952 -22552
rect 21410 -22608 21470 -22548
rect 22922 -22608 22982 -22548
rect 19870 -22738 19930 -22678
rect 20396 -22736 20456 -22676
rect 11724 -23654 11784 -23594
rect 13766 -23654 13826 -23594
rect 15802 -23654 15862 -23594
rect 11220 -23768 11280 -23708
rect 16308 -23764 16368 -23704
rect 10712 -23882 10772 -23822
rect 12742 -23882 12802 -23822
rect 14780 -23882 14840 -23822
rect 16816 -23882 16876 -23822
rect 10556 -23986 10616 -23926
rect 7654 -24988 7714 -24928
rect 7154 -25094 7214 -25034
rect 8168 -25094 8228 -25034
rect 6640 -25204 6700 -25144
rect 5110 -26234 5170 -26174
rect 6132 -26234 6192 -26174
rect 9848 -24882 9908 -24822
rect 9694 -24988 9754 -24928
rect 9200 -25094 9260 -25034
rect 8678 -25204 8738 -25144
rect 7654 -26126 7714 -26066
rect 7146 -26234 7206 -26174
rect 8172 -26234 8232 -26174
rect 10212 -25094 10272 -25034
rect 11726 -24882 11786 -24822
rect 11730 -24988 11790 -24928
rect 11220 -25094 11280 -25034
rect 10716 -25204 10776 -25144
rect 9184 -26234 9244 -26174
rect 10220 -26234 10280 -26174
rect 12238 -25094 12298 -25034
rect 13764 -24882 13824 -24822
rect 13766 -24988 13826 -24928
rect 13264 -25094 13324 -25034
rect 12752 -25204 12812 -25144
rect 11226 -26234 11286 -26174
rect 12240 -26234 12300 -26174
rect 14266 -25094 14326 -25034
rect 16962 -23986 17022 -23926
rect 21910 -22736 21970 -22676
rect 17838 -23882 17898 -23822
rect 18856 -23654 18916 -23594
rect 18858 -23882 18918 -23822
rect 15634 -24882 15694 -24822
rect 15286 -25094 15346 -25034
rect 15800 -24988 15860 -24928
rect 14788 -25204 14848 -25144
rect 13256 -26234 13316 -26174
rect 14264 -26234 14324 -26174
rect 16306 -25094 16366 -25034
rect 19872 -23882 19932 -23822
rect 19872 -23986 19932 -23926
rect 20888 -23654 20948 -23594
rect 23162 -18718 23222 -18658
rect 23400 -18940 23460 -18880
rect 23278 -19042 23338 -18982
rect 23162 -20276 23222 -20216
rect 23158 -21178 23218 -21118
rect 23278 -22404 23338 -22344
rect 23158 -22502 23218 -22442
rect 23034 -23654 23094 -23594
rect 21408 -23764 21468 -23704
rect 22416 -23764 22476 -23704
rect 23526 -20174 23586 -20114
rect 23528 -22608 23588 -22548
rect 23400 -22736 23460 -22676
rect 23762 -16586 23822 -16526
rect 23650 -23764 23710 -23704
rect 20894 -23882 20954 -23822
rect 17840 -24988 17900 -24928
rect 17332 -25094 17392 -25034
rect 18350 -25094 18410 -25034
rect 16820 -25204 16880 -25144
rect 15280 -26234 15340 -26174
rect 16304 -26234 16364 -26174
rect 19870 -24988 19930 -24928
rect 19364 -25094 19424 -25034
rect 18852 -25204 18912 -25144
rect 17834 -26126 17894 -26066
rect 17326 -26234 17386 -26174
rect 18348 -26234 18408 -26174
rect 20378 -25094 20438 -25034
rect 23054 -23986 23114 -23926
rect 21910 -24882 21970 -24822
rect 21910 -24988 21970 -24928
rect 21400 -25094 21460 -25034
rect 20892 -25204 20952 -25144
rect 19366 -26234 19426 -26174
rect 20380 -26234 20440 -26174
rect 23762 -24988 23822 -24928
rect 23054 -26126 23114 -26066
rect 21404 -26234 21464 -26174
rect -8072 -26630 23928 -26476
rect -12216 -27116 -11616 -26816
rect 24216 -27116 24816 -26816
<< metal2 >>
rect 484 4216 1084 4226
rect 484 3906 1084 3916
rect 24116 4216 24716 4226
rect 24116 3906 24716 3916
rect 3998 3834 20878 3866
rect 3998 3620 4061 3834
rect 20846 3620 20878 3834
rect 3998 3600 20878 3620
rect 3998 3598 8352 3600
rect 7986 1918 8046 1924
rect 9068 1918 9128 1924
rect 10026 1918 10086 1924
rect 13090 1918 13150 1924
rect 14108 1918 14168 1924
rect 15132 1918 15192 1924
rect 16144 1918 16204 1924
rect 19202 1918 19262 1924
rect 20214 1918 20274 1924
rect 21232 1918 21292 1924
rect 8046 1858 9068 1918
rect 9128 1858 10026 1918
rect 10086 1858 13090 1918
rect 13150 1858 14108 1918
rect 14168 1858 15132 1918
rect 15192 1858 16144 1918
rect 16204 1858 19202 1918
rect 19262 1858 20214 1918
rect 20274 1858 21232 1918
rect 7986 1852 8046 1858
rect 9068 1852 9128 1858
rect 10026 1852 10086 1858
rect 13090 1852 13150 1858
rect 14108 1852 14168 1858
rect 15132 1852 15192 1858
rect 16144 1852 16204 1858
rect 19202 1852 19262 1858
rect 20214 1852 20274 1858
rect 21232 1852 21292 1858
rect 8512 1672 8572 1678
rect 10548 1672 10608 1678
rect 12586 1674 12646 1680
rect 14616 1674 14676 1680
rect 16658 1676 16718 1682
rect 17668 1676 17728 1682
rect 18690 1676 18750 1682
rect 20726 1676 20786 1682
rect 8572 1612 10548 1672
rect 10608 1614 12586 1672
rect 12646 1614 14616 1674
rect 14676 1616 16658 1674
rect 16718 1616 17668 1676
rect 17728 1616 18690 1676
rect 18750 1616 20726 1676
rect 14676 1614 16856 1616
rect 10608 1612 12768 1614
rect 8512 1606 8572 1612
rect 10548 1606 10608 1612
rect 12586 1608 12646 1612
rect 14616 1608 14676 1614
rect 16658 1610 16718 1614
rect 17668 1610 17728 1616
rect 18690 1610 18750 1616
rect 20726 1610 20786 1616
rect 6330 740 6390 746
rect 7494 740 7554 746
rect 13604 740 13664 746
rect 6390 680 7494 740
rect 7554 680 13604 740
rect 6330 674 6390 680
rect 7494 674 7554 680
rect 13604 674 13664 680
rect 15638 740 15698 746
rect 21746 740 21806 746
rect 22996 740 23056 746
rect 15698 680 21746 740
rect 21806 680 22996 740
rect 15638 674 15698 680
rect 21746 674 21806 680
rect 22996 674 23056 680
rect 9530 636 9590 642
rect 11566 636 11626 642
rect 17672 636 17732 642
rect 19706 636 19766 642
rect 9590 576 11566 636
rect 11626 628 12044 636
rect 12260 628 17672 636
rect 11626 582 17672 628
rect 11626 578 14060 582
rect 11626 576 13034 578
rect 13272 576 14060 578
rect 14276 576 17672 582
rect 17732 576 19706 636
rect 9530 570 9590 576
rect 11566 570 11626 576
rect 17672 570 17732 576
rect 19706 570 19766 576
rect 6200 536 6260 542
rect 7494 536 7554 542
rect 13600 536 13660 542
rect 15636 536 15696 542
rect 6260 476 7494 536
rect 7554 476 13600 536
rect 13660 476 15636 536
rect 6200 470 6260 476
rect 7494 470 7554 476
rect 13600 470 13660 476
rect 15636 470 15696 476
rect 16138 536 16198 542
rect 17158 536 17218 542
rect 18184 536 18244 542
rect 16198 476 17158 536
rect 17218 476 18184 536
rect 16138 470 16198 476
rect 17158 470 17218 476
rect 18184 470 18244 476
rect 18690 532 18750 538
rect 19204 532 19264 538
rect 19708 532 19768 538
rect 20214 532 20274 538
rect 18750 472 19204 532
rect 19264 472 19708 532
rect 19768 472 20214 532
rect 20274 472 20734 532
rect 20794 472 20800 532
rect 18690 466 18750 472
rect 19204 466 19264 472
rect 19708 466 19768 472
rect 20214 466 20274 472
rect 10546 -398 10606 -392
rect 12580 -398 12640 -392
rect 14618 -398 14678 -394
rect 10030 -458 10036 -398
rect 10096 -458 10546 -398
rect 10606 -458 12580 -398
rect 12640 -400 14822 -398
rect 16654 -400 16714 -394
rect 17154 -400 17214 -394
rect 17668 -400 17728 -394
rect 18192 -400 18252 -394
rect 18690 -400 18750 -394
rect 19192 -400 19252 -394
rect 12640 -458 14618 -400
rect 10546 -464 10606 -458
rect 12580 -464 12640 -458
rect 14678 -460 16654 -400
rect 16714 -460 17154 -400
rect 17214 -460 17668 -400
rect 17728 -460 18192 -400
rect 18252 -460 18690 -400
rect 18750 -460 19192 -400
rect 19252 -402 19560 -400
rect 19706 -402 19766 -396
rect 20214 -402 20274 -396
rect 20724 -402 20784 -396
rect 19252 -460 19706 -402
rect 14618 -466 14678 -460
rect 16654 -466 16714 -460
rect 17154 -466 17214 -460
rect 17668 -466 17728 -460
rect 18192 -466 18252 -460
rect 18589 -462 19104 -460
rect 18690 -466 18750 -462
rect 19192 -466 19252 -460
rect 19354 -462 19706 -460
rect 19766 -462 20214 -402
rect 20274 -462 20724 -402
rect 19706 -468 19766 -462
rect 20214 -468 20274 -462
rect 20724 -468 20784 -462
rect 9528 -496 9592 -490
rect 11404 -496 11468 -490
rect 9592 -560 11404 -496
rect 9528 -566 9592 -560
rect 11404 -566 11468 -560
rect 15638 -498 15698 -492
rect 21746 -498 21806 -492
rect 15698 -558 21746 -498
rect 15638 -564 15698 -558
rect 21746 -564 21806 -558
rect 11040 -606 11100 -600
rect 12064 -606 12124 -600
rect 13092 -606 13152 -600
rect 9018 -614 9078 -608
rect 10030 -614 10090 -608
rect 7974 -674 7980 -614
rect 8040 -674 9018 -614
rect 9078 -674 10030 -614
rect 11100 -666 12064 -606
rect 12124 -666 13092 -606
rect 11040 -672 11100 -666
rect 12064 -672 12124 -666
rect 13092 -672 13152 -666
rect 19196 -614 19256 -608
rect 20208 -614 20268 -608
rect 21210 -614 21270 -608
rect 9018 -680 9078 -674
rect 10030 -680 10090 -674
rect 19256 -674 20208 -614
rect 20268 -674 21210 -614
rect 19196 -680 19256 -674
rect 20208 -680 20268 -674
rect 21210 -680 21270 -674
rect 8510 -1536 8570 -1530
rect 10546 -1536 10606 -1530
rect 11068 -1536 11128 -1530
rect 11566 -1536 11626 -1530
rect 12580 -1536 12640 -1530
rect 13040 -1536 13100 -1530
rect 14078 -1536 14084 -1534
rect 8570 -1596 10546 -1536
rect 10606 -1596 11068 -1536
rect 11128 -1596 11566 -1536
rect 11626 -1538 12580 -1536
rect 11626 -1540 12548 -1538
rect 11626 -1596 12040 -1540
rect 8510 -1602 8570 -1596
rect 10546 -1602 10606 -1596
rect 11068 -1602 11128 -1596
rect 11566 -1602 11626 -1596
rect 12034 -1600 12040 -1596
rect 12100 -1596 12548 -1540
rect 12640 -1596 13040 -1536
rect 13100 -1594 14084 -1536
rect 14144 -1536 14150 -1534
rect 14616 -1536 14676 -1530
rect 16122 -1536 16128 -1534
rect 14144 -1594 14616 -1536
rect 13100 -1596 14616 -1594
rect 14676 -1594 16128 -1536
rect 16188 -1536 16194 -1534
rect 16188 -1538 16500 -1536
rect 16654 -1538 16714 -1532
rect 18690 -1538 18750 -1534
rect 16188 -1540 16654 -1538
rect 16714 -1540 18878 -1538
rect 20724 -1540 20784 -1534
rect 16188 -1594 16622 -1540
rect 14676 -1596 16622 -1594
rect 12100 -1600 12106 -1596
rect 12542 -1598 12548 -1596
rect 12608 -1598 12640 -1596
rect 12580 -1602 12640 -1598
rect 13040 -1602 13100 -1596
rect 14616 -1602 14676 -1596
rect 14760 -1598 16086 -1596
rect 16292 -1598 16622 -1596
rect 16714 -1544 17638 -1540
rect 17698 -1542 18690 -1540
rect 16714 -1598 17150 -1544
rect 16616 -1600 16622 -1598
rect 16682 -1600 16714 -1598
rect 16654 -1604 16714 -1600
rect 17144 -1604 17150 -1598
rect 17210 -1598 17638 -1544
rect 17210 -1604 17216 -1598
rect 17632 -1600 17638 -1598
rect 17732 -1544 18690 -1542
rect 17732 -1598 18150 -1544
rect 17666 -1602 17672 -1600
rect 17732 -1602 17738 -1598
rect 18144 -1604 18150 -1598
rect 18210 -1598 18690 -1544
rect 18210 -1604 18216 -1598
rect 18750 -1600 20724 -1540
rect 18690 -1606 18750 -1600
rect 20724 -1606 20784 -1600
rect 4192 -1646 4252 -1642
rect 9526 -1646 9590 -1640
rect 19706 -1646 19770 -1640
rect 4190 -1648 9526 -1646
rect 4190 -1708 4192 -1648
rect 4252 -1708 9526 -1648
rect 4190 -1710 9526 -1708
rect 9590 -1710 19706 -1646
rect 4192 -1714 4252 -1710
rect 9526 -1716 9590 -1710
rect 19706 -1716 19770 -1710
rect 7488 -1784 7552 -1778
rect 7552 -1788 22992 -1784
rect 7552 -1848 13598 -1788
rect 7488 -1854 7552 -1848
rect 13592 -1852 13598 -1848
rect 13662 -1848 22992 -1788
rect 23056 -1848 23062 -1784
rect 13662 -1852 13668 -1848
rect 6330 -1934 6390 -1928
rect 15634 -1930 15698 -1924
rect 6390 -1994 7312 -1934
rect 7372 -1994 15634 -1934
rect 21740 -1934 21800 -1928
rect 15698 -1994 21740 -1934
rect 6330 -2000 6390 -1994
rect 15634 -2000 15698 -1994
rect 21740 -2000 21800 -1994
rect 7428 -2040 7488 -2034
rect 7990 -2040 8050 -2034
rect 9032 -2040 9092 -2034
rect 10032 -2040 10092 -2034
rect 13194 -2040 13254 -2034
rect 14204 -2040 14264 -2034
rect 15146 -2040 15206 -2034
rect 7488 -2100 7990 -2040
rect 8050 -2100 9032 -2040
rect 9092 -2100 10032 -2040
rect 10092 -2100 13194 -2040
rect 13254 -2100 14204 -2040
rect 14264 -2100 15146 -2040
rect 7428 -2106 7488 -2100
rect 7990 -2106 8050 -2100
rect 9032 -2106 9092 -2100
rect 10032 -2106 10092 -2100
rect 13194 -2106 13254 -2100
rect 14204 -2106 14264 -2100
rect 15146 -2106 15206 -2100
rect 7542 -2242 7602 -2236
rect 10720 -2242 10780 -2236
rect 14788 -2242 14848 -2236
rect 18864 -2242 18924 -2236
rect 22060 -2242 22120 -2236
rect 7602 -2302 10720 -2242
rect 10780 -2302 14788 -2242
rect 14848 -2302 18864 -2242
rect 18924 -2302 22060 -2242
rect 7542 -2308 7602 -2302
rect 10720 -2308 10780 -2302
rect 14788 -2308 14848 -2302
rect 18864 -2308 18924 -2302
rect 22060 -2308 22120 -2302
rect 8686 -3178 8746 -3172
rect 10720 -3178 10780 -3172
rect 12762 -3178 12822 -3172
rect 14788 -3178 14848 -3172
rect 16830 -3178 16890 -3172
rect 18866 -3178 18926 -3172
rect 20902 -3178 20962 -3172
rect 8746 -3238 10720 -3178
rect 10780 -3238 12762 -3178
rect 12822 -3238 14788 -3178
rect 14848 -3238 16830 -3178
rect 16890 -3238 18866 -3178
rect 18926 -3238 20902 -3178
rect 8686 -3244 8746 -3238
rect 10720 -3244 10780 -3238
rect 12762 -3244 12822 -3238
rect 14788 -3244 14848 -3238
rect 16830 -3244 16890 -3238
rect 18866 -3244 18926 -3238
rect 20902 -3244 20962 -3238
rect 9190 -3286 9250 -3280
rect 9250 -3346 10212 -3286
rect 10272 -3346 11230 -3286
rect 11290 -3346 12254 -3286
rect 12314 -3346 13268 -3286
rect 13328 -3346 14286 -3286
rect 14346 -3346 15296 -3286
rect 15356 -3346 16318 -3286
rect 16378 -3346 17332 -3286
rect 17392 -3346 18364 -3286
rect 18424 -3346 19374 -3286
rect 19434 -3346 20396 -3286
rect 20456 -3346 20462 -3286
rect 9190 -3352 9250 -3346
rect 8682 -4210 8742 -4204
rect 12762 -4210 12822 -4204
rect 16830 -4210 16890 -4204
rect 20898 -4210 20958 -4204
rect 23290 -4210 23350 -4204
rect 1150 -4270 8682 -4210
rect 8742 -4270 12762 -4210
rect 12822 -4270 16830 -4210
rect 16890 -4270 20898 -4210
rect 20958 -4270 23290 -4210
rect -13992 -10378 -2722 -10122
rect -13992 -10670 -13630 -10378
rect -2866 -10670 -2722 -10378
rect -13992 -10978 -2722 -10670
rect -13992 -11300 -1640 -10978
rect 1150 -11622 1210 -4270
rect 8682 -4276 8742 -4270
rect 12762 -4276 12822 -4270
rect 16830 -4276 16890 -4270
rect 20898 -4276 20958 -4270
rect 23290 -4276 23350 -4270
rect 6686 -4342 6746 -4336
rect 11228 -4342 11234 -4340
rect 6746 -4344 11234 -4342
rect 6746 -4402 9188 -4344
rect 6686 -4408 6746 -4402
rect 9182 -4404 9188 -4402
rect 9248 -4348 11234 -4344
rect 9248 -4402 10202 -4348
rect 9248 -4404 9254 -4402
rect 10196 -4408 10202 -4402
rect 10262 -4400 11234 -4348
rect 11294 -4342 11300 -4340
rect 12226 -4342 12232 -4340
rect 11294 -4400 12232 -4342
rect 12292 -4342 12298 -4340
rect 13270 -4342 13276 -4340
rect 12292 -4400 13276 -4342
rect 13336 -4342 13342 -4340
rect 17326 -4342 17332 -4340
rect 13336 -4344 17332 -4342
rect 13336 -4400 14280 -4344
rect 10262 -4402 14280 -4400
rect 10262 -4408 10268 -4402
rect 14274 -4404 14280 -4402
rect 14340 -4402 15296 -4344
rect 14340 -4404 14346 -4402
rect 15290 -4404 15296 -4402
rect 15356 -4402 16300 -4344
rect 15356 -4404 15362 -4402
rect 16294 -4404 16300 -4402
rect 16360 -4400 17332 -4344
rect 17392 -4342 17398 -4340
rect 22854 -4342 22914 -4336
rect 17392 -4344 22854 -4342
rect 17392 -4400 18348 -4344
rect 16360 -4402 18348 -4400
rect 16360 -4404 16366 -4402
rect 18342 -4404 18348 -4402
rect 18408 -4402 19376 -4344
rect 18408 -4404 18414 -4402
rect 19370 -4404 19376 -4402
rect 19436 -4402 20396 -4344
rect 19436 -4404 19442 -4402
rect 20390 -4404 20396 -4402
rect 20456 -4402 22854 -4344
rect 20456 -4404 20462 -4402
rect 22854 -4408 22914 -4402
rect 14080 -4552 14140 -4546
rect 14140 -4612 15816 -4552
rect 15876 -4612 15882 -4552
rect 21714 -4566 21774 -4562
rect 21712 -4568 23056 -4566
rect 14080 -4618 14140 -4612
rect 21712 -4628 21714 -4568
rect 21774 -4570 23056 -4568
rect 21774 -4628 22996 -4570
rect 21712 -4630 22996 -4628
rect 23056 -4630 23062 -4570
rect 21714 -4634 21774 -4630
rect 15096 -4748 15160 -4742
rect 19160 -4748 19224 -4742
rect 20184 -4748 20248 -4742
rect 21196 -4748 21260 -4742
rect 15160 -4812 19160 -4748
rect 19224 -4812 20184 -4748
rect 20248 -4812 21196 -4748
rect 15096 -4818 15160 -4812
rect 19160 -4818 19224 -4812
rect 20184 -4818 20248 -4812
rect 21196 -4818 21260 -4812
rect 7312 -4870 7372 -4864
rect 8478 -4870 8538 -4864
rect 10514 -4870 10574 -4864
rect 7372 -4930 8478 -4870
rect 8538 -4930 10514 -4870
rect 7312 -4936 7372 -4930
rect 8478 -4936 8538 -4930
rect 10514 -4936 10574 -4930
rect 11022 -4870 11086 -4864
rect 15098 -4870 15162 -4864
rect 11086 -4934 15098 -4870
rect 11022 -4940 11086 -4934
rect 15098 -4940 15162 -4934
rect 18660 -4870 18720 -4864
rect 20694 -4870 20754 -4864
rect 23138 -4870 23198 -4864
rect 18720 -4930 20694 -4870
rect 20754 -4930 23138 -4870
rect 18660 -4936 18720 -4930
rect 20694 -4936 20754 -4930
rect 23138 -4936 23198 -4930
rect 6560 -4952 6620 -4946
rect 6802 -4952 6862 -4946
rect 6620 -5012 6802 -4952
rect 6560 -5018 6620 -5012
rect 6802 -5018 6862 -5012
rect 9496 -5818 9556 -5812
rect 11532 -5818 11592 -5812
rect 9556 -5878 11532 -5818
rect 9496 -5884 9556 -5878
rect 11532 -5884 11592 -5878
rect 11874 -5816 11934 -5810
rect 14588 -5816 14648 -5810
rect 11934 -5876 14588 -5816
rect 11874 -5882 11934 -5876
rect 14588 -5882 14648 -5876
rect 19676 -5818 19736 -5812
rect 21712 -5818 21772 -5812
rect 19736 -5878 21712 -5818
rect 19676 -5884 19736 -5878
rect 3676 -5906 3736 -5900
rect 4698 -5906 4758 -5900
rect 3736 -5966 4698 -5906
rect 3676 -5972 3736 -5966
rect 4698 -5972 4758 -5966
rect 7044 -5916 7104 -5910
rect 19784 -5916 19844 -5878
rect 21712 -5884 21772 -5878
rect 7104 -5976 19844 -5916
rect 7044 -5982 7104 -5976
rect 3784 -6018 3844 -6012
rect 4568 -6018 4628 -6012
rect 3844 -6078 4568 -6018
rect 3784 -6084 3844 -6078
rect 4568 -6084 4628 -6078
rect 7180 -6014 7240 -6008
rect 9496 -6014 9556 -6008
rect 7240 -6074 9496 -6014
rect 7180 -6080 7240 -6074
rect 9496 -6080 9556 -6074
rect 10516 -6012 10576 -6006
rect 15606 -6012 15666 -6006
rect 22978 -6012 23038 -6006
rect 10576 -6072 15606 -6012
rect 15666 -6072 22978 -6012
rect 10516 -6078 10576 -6072
rect 15606 -6078 15666 -6072
rect 22978 -6078 23038 -6072
rect 8482 -6124 8542 -6118
rect 10516 -6124 10576 -6118
rect 8542 -6184 10516 -6124
rect 8482 -6190 8542 -6184
rect 10516 -6190 10576 -6184
rect 13572 -6126 13632 -6120
rect 15606 -6126 15666 -6120
rect 13632 -6186 15606 -6126
rect 13572 -6192 13632 -6186
rect 15606 -6192 15666 -6186
rect 18662 -6126 18722 -6120
rect 20696 -6124 20756 -6120
rect 20628 -6126 20756 -6124
rect 23290 -6126 23350 -6120
rect 18722 -6186 20696 -6126
rect 20756 -6186 23290 -6126
rect 18662 -6192 18722 -6186
rect 20628 -6188 20756 -6186
rect 20696 -6192 20756 -6188
rect 23290 -6192 23350 -6186
rect 2014 -6940 2074 -6934
rect 5208 -6940 5268 -6934
rect 2074 -7000 5208 -6940
rect 2014 -7006 2074 -7000
rect 5208 -7006 5268 -7000
rect 3174 -7050 3234 -7044
rect 6360 -7050 6420 -7044
rect 3234 -7110 6360 -7050
rect 19526 -7060 19586 -7054
rect 3174 -7116 3234 -7110
rect 6360 -7116 6420 -7110
rect 6802 -7074 6862 -7068
rect 13568 -7074 13628 -7068
rect 14588 -7074 14648 -7068
rect 16624 -7074 16684 -7068
rect 6862 -7134 13568 -7074
rect 13628 -7134 14588 -7074
rect 14648 -7134 16624 -7074
rect 19586 -7120 23948 -7060
rect 19526 -7126 19586 -7120
rect 6802 -7140 6862 -7134
rect 13568 -7140 13628 -7134
rect 14588 -7140 14648 -7134
rect 16624 -7140 16684 -7134
rect 19674 -7170 19734 -7164
rect 21714 -7170 21774 -7164
rect 22854 -7170 22914 -7164
rect 6552 -7178 6612 -7172
rect 11534 -7178 11594 -7172
rect 18658 -7178 18718 -7172
rect 6612 -7238 9498 -7178
rect 9558 -7238 11534 -7178
rect 11594 -7238 18658 -7178
rect 19734 -7230 21714 -7170
rect 21774 -7230 22854 -7170
rect 19674 -7236 19734 -7230
rect 21714 -7236 21774 -7230
rect 22854 -7236 22914 -7230
rect 6552 -7244 6612 -7238
rect 11534 -7244 11594 -7238
rect 18658 -7244 18718 -7238
rect 11532 -7280 11592 -7274
rect 20694 -7280 20754 -7274
rect 6798 -7288 6858 -7282
rect 7464 -7288 7524 -7282
rect 6858 -7348 7464 -7288
rect 11592 -7340 20694 -7280
rect 11532 -7346 11592 -7340
rect 20694 -7346 20754 -7340
rect 6798 -7354 6858 -7348
rect 7464 -7354 7524 -7348
rect 9498 -7382 9558 -7376
rect 11532 -7382 11592 -7376
rect 9558 -7442 11532 -7382
rect 9498 -7448 9558 -7442
rect 11532 -7448 11592 -7442
rect 14588 -7380 14648 -7374
rect 15606 -7380 15666 -7374
rect 16622 -7380 16682 -7374
rect 19526 -7380 19586 -7374
rect 14648 -7440 15606 -7380
rect 15666 -7440 16622 -7380
rect 16682 -7440 19526 -7380
rect 14588 -7446 14648 -7440
rect 15606 -7446 15666 -7440
rect 16622 -7446 16682 -7440
rect 19526 -7446 19586 -7440
rect 19678 -7378 19738 -7372
rect 21712 -7378 21772 -7372
rect 22978 -7378 23038 -7372
rect 19738 -7438 21712 -7378
rect 21772 -7438 22978 -7378
rect 23038 -7438 23820 -7378
rect 19678 -7444 19738 -7438
rect 21712 -7444 21772 -7438
rect 22978 -7444 23038 -7438
rect 3690 -7974 3750 -7968
rect 4700 -7974 4760 -7968
rect 1882 -8088 1888 -8028
rect 1948 -8088 1954 -8028
rect 3750 -8034 4700 -7974
rect 3690 -8040 3750 -8034
rect 4700 -8040 4760 -8034
rect 3796 -8074 3856 -8068
rect 4582 -8074 4642 -8068
rect 1396 -9144 1402 -9084
rect 1462 -9144 1468 -9084
rect 1276 -9644 1282 -9584
rect 1342 -9644 1348 -9584
rect 1282 -11494 1342 -9644
rect 1282 -11560 1342 -11554
rect 1402 -11492 1462 -9144
rect 1536 -9320 1542 -9260
rect 1602 -9320 1608 -9260
rect 1542 -11474 1602 -9320
rect 1764 -10142 1770 -10082
rect 1830 -10142 1836 -10082
rect 1770 -11458 1830 -10142
rect 1888 -11358 1948 -8088
rect 3856 -8134 4582 -8074
rect 3796 -8140 3856 -8134
rect 4582 -8140 4642 -8134
rect 11534 -8322 11594 -8316
rect 13336 -8322 13396 -8316
rect 6686 -8330 6746 -8324
rect 8480 -8330 8540 -8324
rect 10516 -8330 10576 -8324
rect 6746 -8390 8480 -8330
rect 8540 -8390 10516 -8330
rect 11594 -8382 13336 -8322
rect 11534 -8388 11594 -8382
rect 13336 -8388 13396 -8382
rect 13570 -8328 13630 -8322
rect 15606 -8328 15666 -8322
rect 13630 -8388 15606 -8328
rect 6686 -8396 6746 -8390
rect 2436 -9494 2442 -9434
rect 2502 -9494 2508 -9434
rect 2330 -9906 2336 -9846
rect 2396 -9906 2402 -9846
rect 2210 -10024 2216 -9964
rect 2276 -10024 2282 -9964
rect 2216 -11348 2276 -10024
rect 2336 -10940 2396 -9906
rect 2319 -10949 2409 -10940
rect 2319 -11048 2409 -11039
rect 1882 -11418 1888 -11358
rect 1948 -11418 1954 -11358
rect 2336 -11356 2396 -11048
rect 2216 -11414 2276 -11408
rect 2330 -11416 2336 -11356
rect 2396 -11416 2402 -11356
rect 2442 -11492 2502 -9494
rect 1770 -11524 1830 -11518
rect 1542 -11540 1602 -11534
rect 2436 -11552 2442 -11492
rect 2502 -11552 2508 -11492
rect 1402 -11558 1462 -11552
rect 1660 -11612 1720 -11606
rect 6914 -11612 6974 -8390
rect 8480 -8396 8540 -8390
rect 10516 -8396 10576 -8390
rect 13570 -8394 13630 -8388
rect 15606 -8394 15666 -8388
rect 18660 -8326 18720 -8320
rect 20696 -8326 20756 -8320
rect 18720 -8386 20696 -8326
rect 18660 -8392 18720 -8386
rect 20696 -8392 20756 -8386
rect 10516 -8438 10576 -8432
rect 15604 -8438 15664 -8432
rect 22854 -8438 22914 -8432
rect 10576 -8498 15604 -8438
rect 15664 -8498 22854 -8438
rect 10516 -8504 10576 -8498
rect 15604 -8504 15664 -8498
rect 22854 -8504 22914 -8498
rect 7312 -8538 7372 -8532
rect 7372 -8598 19896 -8538
rect 7312 -8604 7372 -8598
rect 9494 -8640 9554 -8634
rect 11528 -8640 11588 -8634
rect 9554 -8700 11528 -8640
rect 19682 -8640 19742 -8634
rect 19836 -8640 19896 -8598
rect 21716 -8640 21776 -8634
rect 9494 -8706 9554 -8700
rect 11528 -8706 11588 -8700
rect 11732 -8652 11792 -8646
rect 11792 -8712 15094 -8652
rect 15154 -8712 16110 -8652
rect 16170 -8712 19170 -8652
rect 19230 -8712 19236 -8652
rect 19742 -8700 21716 -8640
rect 19682 -8706 19742 -8700
rect 21716 -8706 21776 -8700
rect 11732 -8718 11792 -8712
rect 7044 -9588 7104 -9582
rect 8476 -9588 8536 -9582
rect 10512 -9588 10572 -9582
rect 7104 -9648 8476 -9588
rect 8536 -9648 10512 -9588
rect 7044 -9654 7104 -9648
rect 8476 -9654 8536 -9648
rect 10512 -9654 10572 -9648
rect 18664 -9588 18724 -9582
rect 20700 -9588 20760 -9582
rect 18724 -9648 20700 -9588
rect 18664 -9654 18724 -9648
rect 7180 -9718 7240 -9712
rect 18794 -9718 18854 -9648
rect 20700 -9654 20760 -9648
rect 7240 -9778 18854 -9718
rect 7180 -9784 7240 -9778
rect 11534 -9858 11594 -9852
rect 23138 -9858 23198 -9852
rect 11594 -9918 23138 -9858
rect 11534 -9924 11594 -9918
rect 1720 -11672 6974 -11612
rect 1660 -11678 1720 -11672
rect 1150 -11688 1210 -11682
rect 13254 -11842 13314 -9918
rect 13254 -11908 13314 -11902
rect 18358 -11842 18418 -9918
rect 22418 -11848 22478 -9918
rect 23138 -9924 23198 -9918
rect 18358 -11908 18418 -11902
rect 22412 -11908 22418 -11848
rect 22478 -11908 22484 -11848
rect -1562 -12220 -1502 -12214
rect 2216 -12220 2276 -12214
rect -1502 -12280 2216 -12220
rect -1562 -12286 -1502 -12280
rect 2216 -12286 2276 -12280
rect -36 -12354 24 -12348
rect 1770 -12354 1830 -12348
rect 24 -12414 1770 -12354
rect -36 -12420 24 -12414
rect 1770 -12420 1830 -12414
rect 2012 -13578 2072 -13572
rect 2072 -13638 3586 -13578
rect 3646 -13638 3652 -13578
rect 2012 -13644 2072 -13638
rect 4600 -13794 4660 -13788
rect 6640 -13794 6700 -13788
rect 8680 -13794 8740 -13788
rect 10710 -13794 10770 -13788
rect 12750 -13794 12810 -13788
rect 14782 -13794 14842 -13788
rect 16822 -13794 16882 -13788
rect 18858 -13794 18918 -13788
rect 20892 -13794 20952 -13788
rect 4660 -13854 6640 -13794
rect 6700 -13854 8680 -13794
rect 8740 -13854 10710 -13794
rect 10770 -13854 12750 -13794
rect 12810 -13854 14782 -13794
rect 14842 -13854 16822 -13794
rect 16882 -13854 18858 -13794
rect 18918 -13854 20892 -13794
rect 4600 -13860 4660 -13854
rect 6640 -13860 6700 -13854
rect 8680 -13860 8740 -13854
rect 10710 -13860 10770 -13854
rect 12750 -13860 12810 -13854
rect 14782 -13860 14842 -13854
rect 16822 -13860 16882 -13854
rect 18858 -13860 18918 -13854
rect 20892 -13860 20952 -13854
rect 2224 -13914 2284 -13908
rect 2568 -13914 2628 -13908
rect 2284 -13974 2568 -13914
rect 2224 -13980 2284 -13974
rect 2568 -13980 2628 -13974
rect 4092 -13920 4152 -13914
rect 12236 -13920 12296 -13914
rect 4152 -13980 5106 -13920
rect 5166 -13980 6128 -13920
rect 6188 -13980 7142 -13920
rect 7202 -13980 8168 -13920
rect 8228 -13980 9180 -13920
rect 9240 -13980 10216 -13920
rect 10276 -13980 11222 -13920
rect 11282 -13980 12236 -13920
rect 12296 -13980 13252 -13920
rect 13312 -13980 14260 -13920
rect 14320 -13980 15276 -13920
rect 15336 -13980 16300 -13920
rect 16360 -13980 17322 -13920
rect 17382 -13980 18344 -13920
rect 18404 -13980 19362 -13920
rect 19422 -13980 20376 -13920
rect 20436 -13980 21400 -13920
rect 21460 -13980 21466 -13920
rect 4092 -13986 4152 -13980
rect 12236 -13986 12296 -13980
rect 2442 -14036 2502 -14030
rect 7656 -14036 7716 -14030
rect 17844 -14036 17904 -14030
rect 21916 -14036 21976 -14030
rect 23048 -14036 23108 -14030
rect 2502 -14096 7656 -14036
rect 7716 -14096 17844 -14036
rect 17904 -14096 21916 -14036
rect 21976 -14096 23048 -14036
rect 2442 -14102 2502 -14096
rect 7656 -14102 7716 -14096
rect 17844 -14102 17904 -14096
rect 21916 -14102 21976 -14096
rect 23048 -14102 23108 -14096
rect 4604 -14958 4664 -14952
rect 6644 -14958 6704 -14952
rect 8676 -14958 8736 -14952
rect 10708 -14958 10768 -14952
rect 12744 -14958 12804 -14952
rect 14780 -14958 14840 -14952
rect 16818 -14958 16878 -14952
rect 18856 -14958 18916 -14952
rect 20892 -14958 20952 -14952
rect 4664 -15018 6644 -14958
rect 6704 -15018 8676 -14958
rect 8736 -15018 10708 -14958
rect 10768 -15018 12744 -14958
rect 12804 -15018 14780 -14958
rect 14840 -15018 16818 -14958
rect 16878 -15018 18856 -14958
rect 18916 -15018 20892 -14958
rect 4604 -15024 4664 -15018
rect 6644 -15024 6704 -15018
rect 8676 -15024 8736 -15018
rect 10708 -15024 10768 -15018
rect 12744 -15024 12804 -15018
rect 14780 -15024 14840 -15018
rect 16818 -15024 16878 -15018
rect 18856 -15024 18916 -15018
rect 20892 -15024 20952 -15018
rect 4096 -15068 4156 -15062
rect 5118 -15068 5178 -15062
rect 6132 -15068 6192 -15062
rect 7146 -15068 7206 -15062
rect 8164 -15068 8224 -15062
rect 9190 -15068 9250 -15062
rect 10210 -15068 10270 -15062
rect 11230 -15068 11290 -15062
rect 12232 -15068 12292 -15062
rect 13258 -15068 13318 -15062
rect 14276 -15068 14336 -15062
rect 15284 -15068 15344 -15062
rect 16296 -15068 16356 -15062
rect 17328 -15068 17388 -15062
rect 18342 -15068 18402 -15062
rect 19360 -15068 19420 -15062
rect 20384 -15068 20444 -15062
rect 21404 -15068 21464 -15062
rect 4156 -15128 5118 -15068
rect 5178 -15128 6132 -15068
rect 6192 -15128 7146 -15068
rect 7206 -15128 8164 -15068
rect 8224 -15128 9190 -15068
rect 9250 -15128 10210 -15068
rect 10270 -15128 11230 -15068
rect 11290 -15128 12232 -15068
rect 12292 -15128 13258 -15068
rect 13318 -15128 14276 -15068
rect 14336 -15128 15284 -15068
rect 15344 -15128 16296 -15068
rect 16356 -15128 17328 -15068
rect 17388 -15128 18342 -15068
rect 18402 -15128 19360 -15068
rect 19420 -15128 20384 -15068
rect 20444 -15128 21404 -15068
rect 4096 -15134 4156 -15128
rect 5118 -15134 5178 -15128
rect 6132 -15134 6192 -15128
rect 7146 -15134 7206 -15128
rect 8164 -15134 8224 -15128
rect 9190 -15134 9250 -15128
rect 10210 -15134 10270 -15128
rect 11230 -15134 11290 -15128
rect 12232 -15134 12292 -15128
rect 13258 -15134 13318 -15128
rect 14276 -15134 14336 -15128
rect 15284 -15134 15344 -15128
rect 16296 -15134 16356 -15128
rect 17328 -15134 17388 -15128
rect 18342 -15134 18402 -15128
rect 19360 -15134 19420 -15128
rect 20384 -15134 20444 -15128
rect 21404 -15134 21464 -15128
rect 2120 -15174 2180 -15168
rect 3586 -15174 3646 -15168
rect 5626 -15174 5686 -15168
rect 7656 -15174 7716 -15168
rect 9696 -15174 9756 -15168
rect 11730 -15174 11790 -15168
rect 13766 -15174 13826 -15168
rect 15802 -15174 15862 -15168
rect 17842 -15174 17902 -15168
rect 19872 -15174 19932 -15168
rect 21912 -15174 21972 -15168
rect 2180 -15234 3586 -15174
rect 3646 -15234 5626 -15174
rect 5686 -15234 7656 -15174
rect 7716 -15234 9696 -15174
rect 9756 -15234 11730 -15174
rect 11790 -15234 13766 -15174
rect 13826 -15234 15802 -15174
rect 15862 -15234 17842 -15174
rect 17902 -15234 19872 -15174
rect 19932 -15234 21912 -15174
rect 2120 -15240 2180 -15234
rect 3586 -15240 3646 -15234
rect 5626 -15240 5686 -15234
rect 7656 -15240 7716 -15234
rect 9696 -15240 9756 -15234
rect 11730 -15240 11790 -15234
rect 13766 -15240 13826 -15234
rect 15802 -15240 15862 -15234
rect 17842 -15240 17902 -15234
rect 19872 -15240 19932 -15234
rect 21912 -15240 21972 -15234
rect 2572 -15280 2632 -15274
rect 3070 -15280 3130 -15274
rect 3582 -15280 3642 -15274
rect 9862 -15280 9922 -15274
rect 11730 -15280 11790 -15274
rect 13768 -15280 13828 -15274
rect 15648 -15280 15708 -15274
rect 1880 -15340 1886 -15280
rect 1946 -15340 2572 -15280
rect 2632 -15340 3070 -15280
rect 3130 -15340 3582 -15280
rect 3642 -15340 9862 -15280
rect 9922 -15340 11730 -15280
rect 11790 -15340 13768 -15280
rect 13828 -15340 15648 -15280
rect 2572 -15346 2632 -15340
rect 3070 -15346 3130 -15340
rect 3582 -15346 3642 -15340
rect 9862 -15346 9922 -15340
rect 11730 -15346 11790 -15340
rect 13768 -15346 13828 -15340
rect 15648 -15346 15708 -15340
rect 19872 -15278 19932 -15272
rect 23048 -15278 23108 -15272
rect 19932 -15338 23048 -15278
rect 19872 -15344 19932 -15338
rect 23048 -15344 23108 -15338
rect 2442 -16170 2502 -16164
rect 5620 -16170 5680 -16164
rect 8676 -16170 8736 -16164
rect 14782 -16170 14842 -16164
rect 19876 -16170 19936 -16164
rect 2502 -16230 5620 -16170
rect 5680 -16230 8676 -16170
rect 8736 -16230 14782 -16170
rect 14842 -16230 19876 -16170
rect 2442 -16236 2502 -16230
rect 5620 -16236 5680 -16230
rect 8676 -16236 8736 -16230
rect 14782 -16236 14842 -16230
rect 19876 -16236 19936 -16230
rect 2012 -16274 2072 -16268
rect 2566 -16274 2626 -16268
rect 4086 -16274 4146 -16268
rect 2072 -16334 2566 -16274
rect 2626 -16334 4086 -16274
rect 2012 -16340 2072 -16334
rect 2566 -16340 2626 -16334
rect 4086 -16340 4146 -16334
rect 4598 -16274 4658 -16268
rect 5622 -16274 5682 -16268
rect 6634 -16274 6694 -16268
rect 7654 -16274 7714 -16268
rect 10712 -16274 10772 -16268
rect 12750 -16274 12810 -16268
rect 15800 -16274 15860 -16268
rect 16818 -16274 16878 -16268
rect 17838 -16274 17898 -16268
rect 18854 -16274 18914 -16268
rect 20890 -16274 20950 -16268
rect 4658 -16334 5622 -16274
rect 5682 -16334 6634 -16274
rect 6694 -16334 7654 -16274
rect 7714 -16334 10712 -16274
rect 10772 -16334 12750 -16274
rect 12810 -16334 15800 -16274
rect 15860 -16334 16818 -16274
rect 16878 -16334 17838 -16274
rect 17898 -16334 18854 -16274
rect 18914 -16334 20890 -16274
rect 4598 -16340 4658 -16334
rect 5622 -16340 5682 -16334
rect 6634 -16340 6694 -16334
rect 7654 -16340 7714 -16334
rect 10712 -16340 10772 -16334
rect 12750 -16340 12810 -16334
rect 15800 -16340 15860 -16334
rect 16818 -16340 16878 -16334
rect 17838 -16340 17898 -16334
rect 18854 -16340 18914 -16334
rect 20890 -16340 20950 -16334
rect 2336 -16396 2396 -16390
rect 9696 -16396 9756 -16390
rect 11730 -16396 11790 -16390
rect 13760 -16396 13820 -16390
rect 23760 -16396 23820 -7438
rect 2396 -16456 9696 -16396
rect 9756 -16456 11730 -16396
rect 11790 -16456 13760 -16396
rect 13820 -16456 23820 -16396
rect 2336 -16462 2396 -16456
rect 9696 -16462 9756 -16456
rect 11730 -16462 11790 -16456
rect 13760 -16462 13820 -16456
rect 2224 -16510 2284 -16504
rect 3072 -16510 3132 -16504
rect 2284 -16570 3072 -16510
rect 2224 -16576 2284 -16570
rect 3072 -16576 3132 -16570
rect 4604 -16508 4664 -16502
rect 6640 -16508 6700 -16502
rect 23034 -16508 23094 -16502
rect 4664 -16568 6640 -16508
rect 6700 -16568 23034 -16508
rect 4604 -16574 4664 -16568
rect 6640 -16574 6700 -16568
rect 23034 -16574 23094 -16568
rect 23162 -16526 23222 -16520
rect 23762 -16526 23822 -16520
rect 23222 -16586 23762 -16526
rect 23162 -16592 23222 -16586
rect 23762 -16592 23822 -16586
rect 22928 -17396 22988 -17390
rect 23888 -17396 23948 -7120
rect 5620 -17414 5680 -17408
rect 7656 -17414 7716 -17408
rect 15800 -17414 15860 -17408
rect 17836 -17414 17896 -17408
rect 21910 -17414 21970 -17408
rect 2448 -17438 2508 -17432
rect 3586 -17438 3646 -17432
rect 2508 -17498 3586 -17438
rect 3646 -17498 4468 -17438
rect 5680 -17474 7656 -17414
rect 7716 -17474 15800 -17414
rect 15860 -17474 17836 -17414
rect 17896 -17474 21910 -17414
rect 22988 -17456 23948 -17396
rect 22928 -17462 22988 -17456
rect 5620 -17480 5680 -17474
rect 7656 -17480 7716 -17474
rect 15800 -17480 15860 -17474
rect 17836 -17480 17896 -17474
rect 21910 -17480 21970 -17474
rect 2448 -17504 2508 -17498
rect 3586 -17504 3646 -17498
rect 2336 -17638 2396 -17632
rect 3584 -17638 3644 -17632
rect 2396 -17698 3584 -17638
rect 4408 -17634 4468 -17498
rect 4602 -17518 4662 -17512
rect 6642 -17518 6702 -17512
rect 8674 -17518 8734 -17512
rect 10708 -17518 10768 -17512
rect 12748 -17518 12808 -17512
rect 14782 -17518 14842 -17512
rect 4662 -17578 6642 -17518
rect 6702 -17578 8674 -17518
rect 8734 -17578 10708 -17518
rect 10768 -17578 12748 -17518
rect 12808 -17578 14782 -17518
rect 4602 -17584 4662 -17578
rect 6642 -17584 6702 -17578
rect 8674 -17584 8734 -17578
rect 10708 -17584 10768 -17578
rect 12748 -17584 12808 -17578
rect 14782 -17584 14842 -17578
rect 14978 -17522 15038 -17516
rect 19870 -17522 19930 -17516
rect 15038 -17582 19870 -17522
rect 23528 -17526 23588 -17520
rect 14978 -17588 15038 -17582
rect 19870 -17588 19930 -17582
rect 20368 -17586 20374 -17526
rect 20434 -17586 23528 -17526
rect 23528 -17592 23588 -17586
rect 5116 -17632 5176 -17626
rect 8674 -17630 8734 -17624
rect 10710 -17630 10770 -17624
rect 12746 -17630 12806 -17624
rect 14782 -17630 14842 -17624
rect 16816 -17630 16876 -17624
rect 18854 -17630 18914 -17624
rect 20894 -17630 20954 -17624
rect 23278 -17630 23338 -17624
rect 4408 -17692 5116 -17634
rect 5176 -17692 6120 -17632
rect 6180 -17692 7132 -17632
rect 7192 -17692 8152 -17632
rect 8212 -17692 8218 -17632
rect 8734 -17690 10710 -17630
rect 10770 -17690 12746 -17630
rect 12806 -17690 14782 -17630
rect 14842 -17690 16816 -17630
rect 16876 -17690 18854 -17630
rect 18914 -17690 20894 -17630
rect 20954 -17690 23278 -17630
rect 4408 -17694 5458 -17692
rect 5116 -17698 5176 -17694
rect 8674 -17696 8734 -17690
rect 10710 -17696 10770 -17690
rect 12746 -17696 12806 -17690
rect 14782 -17696 14842 -17690
rect 16816 -17696 16876 -17690
rect 18854 -17696 18914 -17690
rect 20894 -17696 20954 -17690
rect 23278 -17696 23338 -17690
rect 2336 -17704 2396 -17698
rect 3584 -17704 3644 -17698
rect 1660 -17740 1720 -17734
rect 2230 -17740 2290 -17734
rect 9692 -17740 9752 -17734
rect 11726 -17740 11786 -17734
rect 13766 -17740 13826 -17734
rect 14978 -17740 15038 -17734
rect 1720 -17800 2230 -17740
rect 2290 -17800 9692 -17740
rect 9752 -17800 11726 -17740
rect 11786 -17800 13766 -17740
rect 13826 -17800 14978 -17740
rect 1660 -17806 1720 -17800
rect 2230 -17806 2290 -17800
rect 9692 -17806 9752 -17800
rect 11726 -17806 11786 -17800
rect 13766 -17806 13826 -17800
rect 14978 -17806 15038 -17800
rect 15272 -17738 15332 -17732
rect 15332 -17798 16300 -17738
rect 16360 -17798 16366 -17738
rect 16818 -17744 16878 -17738
rect 18854 -17744 18914 -17738
rect 20892 -17744 20952 -17738
rect 23034 -17744 23094 -17738
rect 15272 -17804 15332 -17798
rect 16878 -17804 18854 -17744
rect 18914 -17804 20892 -17744
rect 20952 -17804 23034 -17744
rect 16818 -17810 16878 -17804
rect 18854 -17810 18914 -17804
rect 20892 -17810 20952 -17804
rect 23034 -17810 23094 -17804
rect 19366 -18658 19426 -18652
rect 3584 -18670 3644 -18664
rect 5622 -18670 5682 -18664
rect 7658 -18670 7718 -18664
rect 9690 -18670 9750 -18664
rect 3644 -18730 5622 -18670
rect 5682 -18730 7658 -18670
rect 7718 -18730 9690 -18670
rect 14266 -18718 14272 -18658
rect 14332 -18718 19366 -18658
rect 19366 -18724 19426 -18718
rect 19504 -18654 19564 -18648
rect 20386 -18654 20446 -18648
rect 21392 -18654 21452 -18648
rect 19564 -18714 20386 -18654
rect 20446 -18714 21392 -18654
rect 19504 -18720 19564 -18714
rect 20386 -18720 20446 -18714
rect 21392 -18720 21452 -18714
rect 21910 -18658 21970 -18652
rect 23162 -18658 23222 -18652
rect 21970 -18718 23162 -18658
rect 21910 -18724 21970 -18718
rect 23162 -18724 23222 -18718
rect 3584 -18736 3644 -18730
rect 5622 -18736 5682 -18730
rect 7658 -18736 7718 -18730
rect 9690 -18736 9750 -18730
rect 4090 -18772 4150 -18766
rect 9182 -18772 9242 -18766
rect 1150 -18822 1210 -18816
rect 4150 -18832 9182 -18772
rect 4090 -18838 4150 -18832
rect 9182 -18838 9242 -18832
rect 13766 -18786 13826 -18780
rect 21910 -18786 21970 -18780
rect 13826 -18846 21910 -18786
rect 13766 -18852 13826 -18846
rect 21910 -18852 21970 -18846
rect -3398 -19748 -3338 -19742
rect 1150 -19748 1210 -18882
rect 2336 -18874 2396 -18868
rect 5620 -18874 5680 -18868
rect 2396 -18934 5620 -18874
rect 2336 -18940 2396 -18934
rect 5620 -18940 5680 -18934
rect 6128 -18880 6188 -18874
rect 7150 -18880 7210 -18874
rect 8164 -18880 8224 -18874
rect 9182 -18880 9242 -18874
rect 10202 -18880 10262 -18874
rect 17314 -18880 17374 -18874
rect 18344 -18880 18404 -18874
rect 19504 -18880 19564 -18874
rect 6188 -18940 7150 -18880
rect 7210 -18940 8164 -18880
rect 8224 -18940 9182 -18880
rect 9242 -18940 10202 -18880
rect 10262 -18940 17314 -18880
rect 17374 -18940 18344 -18880
rect 18404 -18940 19504 -18880
rect 6128 -18946 6188 -18940
rect 7150 -18946 7210 -18940
rect 8164 -18946 8224 -18940
rect 9182 -18946 9242 -18940
rect 10202 -18946 10262 -18940
rect 17314 -18946 17374 -18940
rect 18344 -18946 18404 -18940
rect 19504 -18946 19564 -18940
rect 19872 -18880 19932 -18874
rect 23400 -18880 23460 -18874
rect 19932 -18940 23400 -18880
rect 19872 -18946 19932 -18940
rect 23400 -18946 23460 -18940
rect 4604 -18974 4664 -18968
rect 6638 -18974 6698 -18968
rect 8674 -18974 8734 -18968
rect 4664 -19034 6638 -18974
rect 6698 -19034 8674 -18974
rect 4604 -19040 4664 -19034
rect 6638 -19040 6698 -19034
rect 8674 -19040 8734 -19034
rect 15802 -18984 15862 -18978
rect 19872 -18984 19932 -18978
rect 15862 -19044 19872 -18984
rect 15802 -19050 15862 -19044
rect 19872 -19050 19932 -19044
rect 20888 -18982 20948 -18976
rect 23278 -18982 23338 -18976
rect 20948 -19042 23278 -18982
rect 20888 -19048 20948 -19042
rect 23278 -19048 23338 -19042
rect -3338 -19808 1210 -19748
rect -3398 -19814 -3338 -19808
rect -5428 -19894 -5368 -19888
rect -1368 -19894 -1308 -19888
rect 816 -19894 876 -19888
rect 1282 -19894 1342 -19888
rect 10710 -19892 10770 -19886
rect 12746 -19892 12806 -19886
rect 14782 -19892 14842 -19886
rect 16820 -19892 16880 -19886
rect -9514 -19954 -9508 -19894
rect -9448 -19954 -5428 -19894
rect -5368 -19954 -1368 -19894
rect -1308 -19954 816 -19894
rect 876 -19954 1282 -19894
rect -5428 -19960 -5368 -19954
rect -1368 -19960 -1308 -19954
rect 816 -19960 876 -19954
rect 1282 -19960 1342 -19954
rect 4086 -19898 4146 -19892
rect 4996 -19898 5056 -19892
rect 5998 -19898 6058 -19892
rect 7150 -19898 7210 -19892
rect 8160 -19898 8220 -19892
rect 9166 -19898 9226 -19892
rect 10210 -19898 10270 -19892
rect 4146 -19958 4996 -19898
rect 5056 -19958 5998 -19898
rect 6058 -19958 7150 -19898
rect 7210 -19958 8160 -19898
rect 8220 -19958 9166 -19898
rect 9226 -19958 10210 -19898
rect 10770 -19952 12746 -19892
rect 12806 -19952 14782 -19892
rect 14842 -19952 16820 -19892
rect 10710 -19958 10770 -19952
rect 12746 -19958 12806 -19952
rect 14782 -19958 14842 -19952
rect 16820 -19958 16880 -19952
rect 18856 -19892 18916 -19886
rect 20894 -19892 20954 -19886
rect 18916 -19952 20894 -19892
rect 18856 -19958 18916 -19952
rect 20894 -19958 20954 -19952
rect 4086 -19964 4146 -19958
rect 4996 -19964 5056 -19958
rect 5998 -19964 6058 -19958
rect 7150 -19964 7210 -19958
rect 8160 -19964 8220 -19958
rect 9166 -19964 9226 -19958
rect 10210 -19964 10270 -19958
rect 6638 -20000 6698 -19994
rect 16812 -20000 16872 -19994
rect 18852 -20000 18912 -19994
rect 20890 -20000 20950 -19994
rect -10662 -20022 -10602 -20016
rect -7984 -20022 -7924 -20016
rect -6952 -20022 -6892 -20016
rect -3892 -20022 -3832 -20016
rect -2896 -20022 -2836 -20016
rect 1402 -20022 1462 -20016
rect -10602 -20082 -7984 -20022
rect -7924 -20082 -6952 -20022
rect -6892 -20082 -3892 -20022
rect -3832 -20082 -2896 -20022
rect -2836 -20082 1402 -20022
rect 6698 -20060 16812 -20000
rect 16872 -20060 18852 -20000
rect 18912 -20060 20890 -20000
rect 6638 -20066 6698 -20060
rect 16812 -20066 16872 -20060
rect 18852 -20066 18912 -20060
rect 20890 -20066 20950 -20060
rect -10662 -20088 -10602 -20082
rect -7984 -20088 -7924 -20082
rect -6952 -20088 -6892 -20082
rect -3892 -20088 -3832 -20082
rect -2896 -20088 -2836 -20082
rect 1402 -20088 1462 -20082
rect 4086 -20114 4146 -20108
rect 6138 -20114 6198 -20108
rect 9164 -20114 9224 -20108
rect 10204 -20114 10264 -20108
rect 11218 -20114 11278 -20108
rect 12226 -20114 12286 -20108
rect 13270 -20114 13330 -20108
rect 14260 -20114 14320 -20108
rect 15278 -20114 15338 -20108
rect 16312 -20114 16372 -20108
rect 19344 -20114 19404 -20108
rect 20382 -20114 20442 -20108
rect 21408 -20114 21468 -20108
rect 4146 -20174 5124 -20114
rect 5184 -20174 6138 -20114
rect 6198 -20174 9164 -20114
rect 9224 -20174 10204 -20114
rect 10264 -20174 11218 -20114
rect 11278 -20174 12226 -20114
rect 12286 -20174 13270 -20114
rect 13330 -20174 14260 -20114
rect 14320 -20174 15278 -20114
rect 15338 -20174 16312 -20114
rect 16372 -20174 19344 -20114
rect 19404 -20174 20382 -20114
rect 20442 -20174 21408 -20114
rect 21468 -20174 23526 -20114
rect 23586 -20174 23592 -20114
rect 4086 -20180 4146 -20174
rect 6138 -20180 6198 -20174
rect 9164 -20180 9224 -20174
rect 10204 -20180 10264 -20174
rect 11218 -20180 11278 -20174
rect 12226 -20180 12286 -20174
rect 13270 -20180 13330 -20174
rect 14260 -20180 14320 -20174
rect 15278 -20180 15338 -20174
rect 16312 -20180 16372 -20174
rect 19344 -20180 19404 -20174
rect 20382 -20180 20442 -20174
rect 21408 -20180 21468 -20174
rect 9688 -20218 9748 -20212
rect 11730 -20218 11790 -20212
rect 13768 -20218 13828 -20212
rect 15802 -20218 15862 -20212
rect 17836 -20216 17896 -20210
rect 19870 -20216 19930 -20210
rect 21912 -20216 21972 -20210
rect 23162 -20216 23222 -20210
rect 2444 -20278 2450 -20218
rect 2510 -20278 9688 -20218
rect 9748 -20278 11730 -20218
rect 11790 -20278 13768 -20218
rect 13828 -20278 15802 -20218
rect 9688 -20284 9748 -20278
rect 11730 -20284 11790 -20278
rect 13768 -20284 13828 -20278
rect 15802 -20284 15862 -20278
rect 16314 -20222 16374 -20216
rect 17336 -20222 17396 -20216
rect 16374 -20282 17336 -20222
rect 17896 -20276 19870 -20216
rect 19930 -20276 21912 -20216
rect 21972 -20276 23162 -20216
rect 17836 -20282 17896 -20276
rect 19870 -20282 19930 -20276
rect 21912 -20282 21972 -20276
rect 23162 -20282 23222 -20276
rect 16314 -20288 16374 -20282
rect 17336 -20288 17396 -20282
rect -9004 -20984 -8944 -20978
rect -7980 -20984 -7920 -20978
rect -6948 -20984 -6888 -20978
rect -5948 -20984 -5888 -20978
rect -4928 -20984 -4868 -20978
rect -3908 -20984 -3848 -20978
rect -1884 -20984 -1824 -20978
rect 936 -20984 996 -20978
rect 1542 -20984 1602 -20978
rect -8944 -21044 -7980 -20984
rect -7920 -21044 -6948 -20984
rect -6888 -21044 -5948 -20984
rect -5888 -21044 -4928 -20984
rect -4868 -21044 -3908 -20984
rect -3848 -21044 -2898 -20984
rect -2838 -21044 -1884 -20984
rect -1824 -21044 -866 -20984
rect -806 -21044 936 -20984
rect 996 -21044 1542 -20984
rect -9004 -21050 -8944 -21044
rect -7980 -21050 -7920 -21044
rect -6948 -21050 -6888 -21044
rect -5948 -21050 -5888 -21044
rect -4928 -21050 -4868 -21044
rect -3908 -21050 -3848 -21044
rect -1884 -21050 -1824 -21044
rect 936 -21050 996 -21044
rect 1542 -21050 1602 -21044
rect -9504 -21088 -9444 -21082
rect -7468 -21088 -7408 -21082
rect -5432 -21088 -5372 -21082
rect -3398 -21088 -3338 -21082
rect -1362 -21088 -1302 -21082
rect -9444 -21148 -7468 -21088
rect -7408 -21148 -5432 -21088
rect -5372 -21148 -3398 -21088
rect -3338 -21148 -1362 -21088
rect 8678 -21120 8738 -21114
rect 12746 -21120 12806 -21114
rect 14780 -21120 14840 -21114
rect -9504 -21154 -9444 -21148
rect -7468 -21154 -7408 -21148
rect -5432 -21154 -5372 -21148
rect -3398 -21154 -3338 -21148
rect -1362 -21154 -1302 -21148
rect 4084 -21126 4144 -21120
rect 5092 -21126 5152 -21120
rect 6106 -21126 6166 -21120
rect 7144 -21126 7204 -21120
rect 8162 -21126 8222 -21120
rect 4144 -21186 5092 -21126
rect 5152 -21186 6106 -21126
rect 6166 -21186 7144 -21126
rect 7204 -21186 8162 -21126
rect 8738 -21180 10714 -21120
rect 10774 -21180 12746 -21120
rect 12806 -21180 14780 -21120
rect 8678 -21186 8738 -21180
rect 12746 -21186 12806 -21180
rect 14780 -21186 14840 -21180
rect 15802 -21118 15862 -21112
rect 16156 -21118 16216 -21112
rect 15862 -21178 16156 -21118
rect 15802 -21184 15862 -21178
rect 16156 -21184 16216 -21178
rect 19874 -21118 19934 -21112
rect 23158 -21118 23218 -21112
rect 19934 -21178 23158 -21118
rect 19874 -21184 19934 -21178
rect 23158 -21184 23218 -21178
rect -4418 -21192 -4358 -21186
rect 2120 -21192 2180 -21186
rect 4084 -21192 4144 -21186
rect 5092 -21192 5152 -21186
rect 6106 -21192 6166 -21186
rect 7144 -21192 7204 -21186
rect 8162 -21192 8222 -21186
rect -8492 -21252 -8486 -21192
rect -8426 -21252 -6450 -21192
rect -6390 -21252 -4418 -21192
rect -4358 -21252 -2384 -21192
rect -2324 -21252 -340 -21192
rect -280 -21252 2120 -21192
rect -4418 -21258 -4358 -21252
rect 2120 -21258 2180 -21252
rect 2230 -21230 2290 -21224
rect 3586 -21230 3646 -21224
rect 11730 -21230 11790 -21224
rect 13766 -21230 13826 -21224
rect 15798 -21230 15858 -21224
rect 2290 -21290 3586 -21230
rect 3646 -21290 11730 -21230
rect 11790 -21290 13766 -21230
rect 13826 -21290 15798 -21230
rect 2230 -21296 2290 -21290
rect 3586 -21296 3646 -21290
rect 11730 -21296 11790 -21290
rect 13766 -21296 13826 -21290
rect 15798 -21296 15858 -21290
rect 15308 -21328 15368 -21322
rect 16346 -21328 16406 -21322
rect 17322 -21328 17382 -21322
rect 18338 -21328 18398 -21322
rect 20364 -21328 20424 -21322
rect 21394 -21328 21454 -21322
rect 1888 -21342 1948 -21336
rect 4602 -21342 4662 -21336
rect 6640 -21342 6700 -21336
rect 10712 -21342 10772 -21336
rect 1948 -21402 4602 -21342
rect 4662 -21402 6640 -21342
rect 6700 -21402 10712 -21342
rect 15368 -21388 16346 -21328
rect 16406 -21388 17322 -21328
rect 17382 -21388 18338 -21328
rect 18398 -21388 20364 -21328
rect 20424 -21388 21394 -21328
rect 15308 -21394 15368 -21388
rect 16346 -21394 16406 -21388
rect 17322 -21394 17382 -21388
rect 18338 -21394 18398 -21388
rect 20364 -21394 20424 -21388
rect 21394 -21394 21454 -21388
rect 1888 -21408 1948 -21402
rect 4602 -21408 4662 -21402
rect 6640 -21408 6700 -21402
rect 10712 -21408 10772 -21402
rect 3582 -21440 3642 -21434
rect 5620 -21440 5680 -21434
rect 7660 -21440 7720 -21434
rect 9696 -21440 9756 -21434
rect 15800 -21440 15860 -21434
rect 16150 -21440 16156 -21436
rect 3642 -21500 5620 -21440
rect 5680 -21500 7660 -21440
rect 7720 -21500 9696 -21440
rect 9756 -21496 16156 -21440
rect 16216 -21440 16222 -21436
rect 17836 -21440 17896 -21434
rect 19872 -21440 19932 -21434
rect 21908 -21440 21968 -21434
rect 16216 -21496 17836 -21440
rect 9756 -21500 17836 -21496
rect 17896 -21500 19872 -21440
rect 19932 -21500 21908 -21440
rect 3582 -21506 3642 -21500
rect 5620 -21506 5680 -21500
rect 7660 -21506 7720 -21500
rect 9696 -21506 9756 -21500
rect 15800 -21506 15860 -21500
rect 17836 -21506 17896 -21500
rect 19872 -21506 19932 -21500
rect 21908 -21506 21968 -21500
rect -7474 -22134 -7414 -22128
rect -3398 -22134 -3338 -22128
rect 816 -22134 876 -22128
rect -7414 -22194 -3398 -22134
rect -3338 -22194 816 -22134
rect -7474 -22200 -7414 -22194
rect -3398 -22200 -3338 -22194
rect 816 -22200 876 -22194
rect -10662 -22254 -10602 -22248
rect -9012 -22254 -8952 -22248
rect -5942 -22254 -5882 -22248
rect -4934 -22254 -4874 -22248
rect -1872 -22254 -1812 -22248
rect -846 -22254 -786 -22248
rect -10602 -22314 -9012 -22254
rect -8952 -22314 -5942 -22254
rect -5882 -22314 -4934 -22254
rect -4874 -22314 -1872 -22254
rect -1812 -22314 -846 -22254
rect -10662 -22320 -10602 -22314
rect -9012 -22320 -8952 -22314
rect -5942 -22320 -5882 -22314
rect -4934 -22320 -4874 -22314
rect -1872 -22320 -1812 -22314
rect -846 -22320 -786 -22314
rect 10708 -22344 10768 -22338
rect 12750 -22344 12810 -22338
rect 14782 -22344 14842 -22338
rect 16822 -22344 16882 -22338
rect 23278 -22344 23338 -22338
rect 4602 -22364 4662 -22358
rect 6638 -22364 6698 -22358
rect 8676 -22364 8736 -22358
rect 4662 -22424 6638 -22364
rect 6698 -22424 8676 -22364
rect 10532 -22404 10538 -22344
rect 10598 -22404 10708 -22344
rect 10768 -22404 12750 -22344
rect 12810 -22404 14782 -22344
rect 14842 -22404 16822 -22344
rect 16882 -22404 23278 -22344
rect 10708 -22410 10768 -22404
rect 12750 -22410 12810 -22404
rect 14782 -22410 14842 -22404
rect 16822 -22410 16882 -22404
rect 23278 -22410 23338 -22404
rect 4602 -22430 4662 -22424
rect 6638 -22430 6698 -22424
rect 8676 -22430 8736 -22424
rect 15800 -22442 15860 -22436
rect 21906 -22442 21966 -22436
rect 23158 -22442 23218 -22436
rect 2448 -22462 2508 -22456
rect 5620 -22462 5680 -22456
rect 2508 -22522 5620 -22462
rect 2448 -22528 2508 -22522
rect 5620 -22528 5680 -22522
rect 7144 -22462 7204 -22456
rect 10192 -22462 10252 -22456
rect 7204 -22522 8166 -22462
rect 8226 -22522 9188 -22462
rect 9248 -22522 10192 -22462
rect 15860 -22502 21906 -22442
rect 21966 -22502 23158 -22442
rect 15800 -22508 15860 -22502
rect 21906 -22508 21966 -22502
rect 23158 -22508 23218 -22502
rect 7144 -22528 7204 -22522
rect 10192 -22528 10252 -22522
rect 10714 -22552 10774 -22546
rect 12742 -22552 12802 -22546
rect 14786 -22552 14846 -22546
rect 16814 -22552 16874 -22546
rect 18852 -22552 18912 -22546
rect 20892 -22552 20952 -22546
rect 4606 -22558 4666 -22552
rect 6642 -22558 6702 -22552
rect 8670 -22558 8730 -22552
rect 10538 -22558 10598 -22552
rect 4666 -22618 6642 -22558
rect 6702 -22618 8670 -22558
rect 8730 -22618 10538 -22558
rect 10774 -22612 12742 -22552
rect 12802 -22612 14786 -22552
rect 14846 -22612 16814 -22552
rect 16874 -22612 18852 -22552
rect 18912 -22612 20892 -22552
rect 10714 -22618 10774 -22612
rect 12742 -22618 12802 -22612
rect 14786 -22618 14846 -22612
rect 16814 -22618 16874 -22612
rect 18852 -22618 18912 -22612
rect 20892 -22618 20952 -22612
rect 21410 -22548 21470 -22542
rect 22922 -22548 22982 -22542
rect 23528 -22548 23588 -22542
rect 21470 -22608 22922 -22548
rect 22982 -22608 23528 -22548
rect 21410 -22614 21470 -22608
rect 22922 -22614 22982 -22608
rect 23528 -22614 23588 -22608
rect 4606 -22624 4666 -22618
rect 6642 -22624 6702 -22618
rect 8670 -22624 8730 -22618
rect 10538 -22624 10598 -22618
rect 3588 -22678 3648 -22672
rect 7656 -22678 7716 -22672
rect 9690 -22678 9750 -22672
rect 17840 -22678 17900 -22672
rect 19870 -22678 19930 -22672
rect 21910 -22676 21970 -22670
rect 23400 -22676 23460 -22670
rect 3648 -22738 7656 -22678
rect 7716 -22738 9690 -22678
rect 9750 -22738 17840 -22678
rect 17900 -22738 19870 -22678
rect 20390 -22736 20396 -22676
rect 20456 -22736 21910 -22676
rect 21970 -22736 23400 -22676
rect 3588 -22744 3648 -22738
rect 7656 -22744 7716 -22738
rect 9690 -22744 9750 -22738
rect 17840 -22744 17900 -22738
rect 19870 -22744 19930 -22738
rect 21910 -22742 21970 -22736
rect 23400 -22742 23460 -22736
rect -340 -23198 -280 -23192
rect -8492 -23258 -8486 -23198
rect -8426 -23258 -6450 -23198
rect -6390 -23258 -4418 -23198
rect -4358 -23258 -2384 -23198
rect -2324 -23258 -340 -23198
rect -340 -23264 -280 -23258
rect -9500 -23306 -9440 -23300
rect -7464 -23306 -7404 -23300
rect -5428 -23306 -5368 -23300
rect -3394 -23306 -3334 -23300
rect -1358 -23306 -1298 -23300
rect -9440 -23366 -7464 -23306
rect -7404 -23366 -5428 -23306
rect -5368 -23366 -3394 -23306
rect -3334 -23366 -1358 -23306
rect -9500 -23372 -9440 -23366
rect -7464 -23372 -7404 -23366
rect -5428 -23372 -5368 -23366
rect -3394 -23372 -3334 -23366
rect -1358 -23372 -1298 -23366
rect -9006 -23418 -8946 -23412
rect -7982 -23418 -7922 -23412
rect -6950 -23418 -6890 -23412
rect -5950 -23418 -5890 -23412
rect -4930 -23418 -4870 -23412
rect -3910 -23418 -3850 -23412
rect -1886 -23418 -1826 -23412
rect 936 -23418 996 -23412
rect -8946 -23478 -7982 -23418
rect -7922 -23478 -6950 -23418
rect -6890 -23478 -5950 -23418
rect -5890 -23478 -4930 -23418
rect -4870 -23478 -3910 -23418
rect -3850 -23478 -2900 -23418
rect -2840 -23478 -1886 -23418
rect -1826 -23478 -868 -23418
rect -808 -23478 936 -23418
rect -9006 -23484 -8946 -23478
rect -7982 -23484 -7922 -23478
rect -6950 -23484 -6890 -23478
rect -5950 -23484 -5890 -23478
rect -4930 -23484 -4870 -23478
rect -3910 -23484 -3850 -23478
rect -1886 -23484 -1826 -23478
rect 936 -23484 996 -23478
rect 2336 -23594 2396 -23588
rect 11724 -23594 11784 -23588
rect 13766 -23594 13826 -23588
rect 15802 -23594 15862 -23588
rect 2396 -23654 11724 -23594
rect 11784 -23654 13766 -23594
rect 13826 -23654 15802 -23594
rect 2336 -23660 2396 -23654
rect 11724 -23660 11784 -23654
rect 13766 -23660 13826 -23654
rect 15802 -23660 15862 -23654
rect 18856 -23594 18916 -23588
rect 20888 -23594 20948 -23588
rect 23034 -23594 23094 -23588
rect 18916 -23654 20888 -23594
rect 20948 -23654 23034 -23594
rect 18856 -23660 18916 -23654
rect 20888 -23660 20948 -23654
rect 23034 -23660 23094 -23654
rect 6140 -23708 6200 -23702
rect 11220 -23708 11280 -23702
rect 2230 -23720 2290 -23714
rect 5620 -23720 5680 -23714
rect 2290 -23780 5620 -23720
rect 6200 -23768 11220 -23708
rect 6140 -23774 6200 -23768
rect 11220 -23774 11280 -23768
rect 16308 -23704 16368 -23698
rect 21408 -23704 21468 -23698
rect 16368 -23764 21408 -23704
rect 16308 -23770 16368 -23764
rect 21408 -23770 21468 -23764
rect 22416 -23704 22476 -23698
rect 23650 -23704 23710 -23698
rect 22476 -23764 23650 -23704
rect 22416 -23770 22476 -23764
rect 23650 -23770 23710 -23764
rect 2230 -23786 2290 -23780
rect 5620 -23786 5680 -23780
rect 4602 -23822 4662 -23816
rect 6638 -23822 6698 -23816
rect 7658 -23822 7718 -23816
rect 8674 -23822 8734 -23816
rect 9694 -23822 9754 -23816
rect 10712 -23822 10772 -23816
rect 12742 -23822 12802 -23816
rect 14780 -23822 14840 -23816
rect 16816 -23822 16876 -23816
rect 17838 -23822 17898 -23816
rect 18858 -23822 18918 -23816
rect 19872 -23822 19932 -23816
rect 20894 -23822 20954 -23816
rect 4662 -23882 6638 -23822
rect 6698 -23882 7658 -23822
rect 7718 -23882 8674 -23822
rect 8734 -23882 9694 -23822
rect 9754 -23882 10712 -23822
rect 10772 -23882 12742 -23822
rect 12802 -23882 14780 -23822
rect 14840 -23882 16816 -23822
rect 16876 -23882 17838 -23822
rect 17898 -23882 18858 -23822
rect 18918 -23882 19872 -23822
rect 19932 -23882 20894 -23822
rect 4602 -23888 4662 -23882
rect 6638 -23888 6698 -23882
rect 7658 -23888 7718 -23882
rect 8674 -23888 8734 -23882
rect 9694 -23888 9754 -23882
rect 10712 -23888 10772 -23882
rect 12742 -23888 12802 -23882
rect 14780 -23888 14840 -23882
rect 16816 -23888 16876 -23882
rect 17838 -23888 17898 -23882
rect 18858 -23888 18918 -23882
rect 19872 -23888 19932 -23882
rect 20894 -23888 20954 -23882
rect 5620 -23926 5680 -23920
rect 10556 -23926 10616 -23920
rect 16962 -23926 17022 -23920
rect 19872 -23926 19932 -23920
rect 23054 -23926 23114 -23920
rect 5680 -23986 10556 -23926
rect 10616 -23986 16962 -23926
rect 17022 -23986 19872 -23926
rect 19932 -23986 23054 -23926
rect 5620 -23992 5680 -23986
rect 10556 -23992 10616 -23986
rect 16962 -23992 17022 -23986
rect 19872 -23992 19932 -23986
rect 23054 -23992 23114 -23986
rect -10662 -24380 -10602 -24374
rect -7992 -24380 -7932 -24374
rect -6960 -24380 -6900 -24374
rect -3900 -24380 -3840 -24374
rect -2904 -24380 -2844 -24374
rect -10602 -24440 -7992 -24380
rect -7932 -24440 -6960 -24380
rect -6900 -24440 -3900 -24380
rect -3840 -24440 -2904 -24380
rect -10662 -24446 -10602 -24440
rect -7992 -24446 -7932 -24440
rect -6960 -24446 -6900 -24440
rect -3900 -24446 -3840 -24440
rect -2904 -24446 -2844 -24440
rect -5426 -24510 -5366 -24504
rect -1366 -24510 -1306 -24504
rect 816 -24510 876 -24504
rect -9512 -24570 -9506 -24510
rect -9446 -24570 -5426 -24510
rect -5366 -24570 -1366 -24510
rect -1306 -24570 816 -24510
rect -5426 -24576 -5366 -24570
rect -1366 -24576 -1306 -24570
rect 816 -24576 876 -24570
rect 2448 -24824 2508 -24818
rect 5618 -24824 5678 -24818
rect 2508 -24884 5618 -24824
rect 2448 -24890 2508 -24884
rect 5618 -24890 5678 -24884
rect 9848 -24822 9908 -24816
rect 11726 -24822 11786 -24816
rect 13764 -24822 13824 -24816
rect 15634 -24822 15694 -24816
rect 21910 -24822 21970 -24816
rect 9908 -24882 11726 -24822
rect 11786 -24882 13764 -24822
rect 13824 -24882 15634 -24822
rect 15694 -24882 21910 -24822
rect 9848 -24888 9908 -24882
rect 11726 -24888 11786 -24882
rect 13764 -24888 13824 -24882
rect 15634 -24888 15694 -24882
rect 21910 -24888 21970 -24882
rect 2120 -24928 2180 -24922
rect 3584 -24928 3644 -24922
rect 5624 -24928 5684 -24922
rect 7654 -24928 7714 -24922
rect 9694 -24928 9754 -24922
rect 11730 -24928 11790 -24922
rect 13766 -24928 13826 -24922
rect 15800 -24928 15860 -24922
rect 17840 -24928 17900 -24922
rect 19870 -24928 19930 -24922
rect 21910 -24928 21970 -24922
rect 23762 -24928 23822 -24922
rect 2180 -24988 3584 -24928
rect 3644 -24988 5624 -24928
rect 5684 -24988 7654 -24928
rect 7714 -24988 9694 -24928
rect 9754 -24988 11730 -24928
rect 11790 -24988 13766 -24928
rect 13826 -24988 15800 -24928
rect 15860 -24988 17840 -24928
rect 17900 -24988 19870 -24928
rect 19930 -24988 21910 -24928
rect 21970 -24988 23762 -24928
rect 2120 -24994 2180 -24988
rect 3584 -24994 3644 -24988
rect 5624 -24994 5684 -24988
rect 7654 -24994 7714 -24988
rect 9694 -24994 9754 -24988
rect 11730 -24994 11790 -24988
rect 13766 -24994 13826 -24988
rect 15800 -24994 15860 -24988
rect 17840 -24994 17900 -24988
rect 19870 -24994 19930 -24988
rect 21910 -24994 21970 -24988
rect 23762 -24994 23822 -24988
rect 4092 -25034 4152 -25028
rect 5112 -25034 5172 -25028
rect 6136 -25034 6196 -25028
rect 7154 -25034 7214 -25028
rect 8168 -25034 8228 -25028
rect 9200 -25034 9260 -25028
rect 10212 -25034 10272 -25028
rect 11220 -25034 11280 -25028
rect 12238 -25034 12298 -25028
rect 13264 -25034 13324 -25028
rect 14266 -25034 14326 -25028
rect 15286 -25034 15346 -25028
rect 16306 -25034 16366 -25028
rect 17332 -25034 17392 -25028
rect 18350 -25034 18410 -25028
rect 19364 -25034 19424 -25028
rect 20378 -25034 20438 -25028
rect 21400 -25034 21460 -25028
rect 4152 -25094 5112 -25034
rect 5172 -25094 6136 -25034
rect 6196 -25094 7154 -25034
rect 7214 -25094 8168 -25034
rect 8228 -25094 9200 -25034
rect 9260 -25094 10212 -25034
rect 10272 -25094 11220 -25034
rect 11280 -25094 12238 -25034
rect 12298 -25094 13264 -25034
rect 13324 -25094 14266 -25034
rect 14326 -25094 15286 -25034
rect 15346 -25094 16306 -25034
rect 16366 -25094 17332 -25034
rect 17392 -25094 18350 -25034
rect 18410 -25094 19364 -25034
rect 19424 -25094 20378 -25034
rect 20438 -25094 21400 -25034
rect 4092 -25100 4152 -25094
rect 5112 -25100 5172 -25094
rect 6136 -25100 6196 -25094
rect 7154 -25100 7214 -25094
rect 8168 -25100 8228 -25094
rect 9200 -25100 9260 -25094
rect 10212 -25100 10272 -25094
rect 11220 -25100 11280 -25094
rect 12238 -25100 12298 -25094
rect 13264 -25100 13324 -25094
rect 14266 -25100 14326 -25094
rect 15286 -25100 15346 -25094
rect 16306 -25100 16366 -25094
rect 17332 -25100 17392 -25094
rect 18350 -25100 18410 -25094
rect 19364 -25100 19424 -25094
rect 20378 -25100 20438 -25094
rect 21400 -25100 21460 -25094
rect 4604 -25144 4664 -25138
rect 6640 -25144 6700 -25138
rect 8678 -25144 8738 -25138
rect 10716 -25144 10776 -25138
rect 12752 -25144 12812 -25138
rect 14788 -25144 14848 -25138
rect 16820 -25144 16880 -25138
rect 18852 -25144 18912 -25138
rect 20892 -25144 20952 -25138
rect 4664 -25204 6640 -25144
rect 6700 -25204 8678 -25144
rect 8738 -25204 10716 -25144
rect 10776 -25204 12752 -25144
rect 12812 -25204 14788 -25144
rect 14848 -25204 16820 -25144
rect 16880 -25204 18852 -25144
rect 18912 -25204 20892 -25144
rect 4604 -25210 4664 -25204
rect 6640 -25210 6700 -25204
rect 8678 -25210 8738 -25204
rect 10716 -25210 10776 -25204
rect 12752 -25210 12812 -25204
rect 14788 -25210 14848 -25204
rect 16820 -25210 16880 -25204
rect 18852 -25210 18912 -25204
rect 20892 -25210 20952 -25204
rect -8028 -25876 -7968 -25870
rect -5990 -25876 -5930 -25870
rect -3954 -25876 -3894 -25870
rect -1918 -25876 -1858 -25870
rect -7968 -25936 -5990 -25876
rect -5930 -25936 -3954 -25876
rect -3894 -25936 -1918 -25876
rect -8028 -25942 -7968 -25936
rect -5990 -25942 -5930 -25936
rect -3954 -25942 -3894 -25936
rect -1918 -25942 -1858 -25936
rect -7010 -25988 -6950 -25982
rect -2936 -25988 -2876 -25982
rect 1070 -25988 1130 -25982
rect -6950 -26048 -2936 -25988
rect -2876 -26048 1070 -25988
rect -7010 -26054 -6950 -26048
rect -2936 -26054 -2876 -26048
rect 1070 -26054 1130 -26048
rect 2448 -26066 2508 -26060
rect 3584 -26066 3644 -26060
rect 7654 -26066 7714 -26060
rect 17834 -26066 17894 -26060
rect 23054 -26066 23114 -26060
rect 2508 -26126 3584 -26066
rect 3644 -26126 7654 -26066
rect 7714 -26126 17834 -26066
rect 17894 -26126 23054 -26066
rect 2448 -26132 2508 -26126
rect 3584 -26132 3644 -26126
rect 7654 -26132 7714 -26126
rect 17834 -26132 17894 -26126
rect 23054 -26132 23114 -26126
rect 4096 -26174 4156 -26168
rect 12240 -26174 12300 -26168
rect 4156 -26234 5110 -26174
rect 5170 -26234 6132 -26174
rect 6192 -26234 7146 -26174
rect 7206 -26234 8172 -26174
rect 8232 -26234 9184 -26174
rect 9244 -26234 10220 -26174
rect 10280 -26234 11226 -26174
rect 11286 -26234 12240 -26174
rect 12300 -26234 13256 -26174
rect 13316 -26234 14264 -26174
rect 14324 -26234 15280 -26174
rect 15340 -26234 16304 -26174
rect 16364 -26234 17326 -26174
rect 17386 -26234 18348 -26174
rect 18408 -26234 19366 -26174
rect 19426 -26234 20380 -26174
rect 20440 -26234 21404 -26174
rect 21464 -26234 21470 -26174
rect 4096 -26240 4156 -26234
rect 12240 -26240 12300 -26234
rect -8118 -26476 23968 -26430
rect -8118 -26630 -8072 -26476
rect 23928 -26630 23968 -26476
rect -8118 -26676 23968 -26630
rect -12216 -26816 -11616 -26806
rect -12216 -27126 -11616 -27116
rect 24216 -26816 24816 -26806
rect 24216 -27126 24816 -27116
<< via2 >>
rect 484 3916 1084 4216
rect 24116 3916 24716 4216
rect 4061 3620 20846 3834
rect -13630 -10670 -2868 -10378
rect 2319 -11039 2409 -10949
rect -8072 -26630 23928 -26476
rect -12216 -27116 -11616 -26816
rect 24216 -27116 24816 -26816
<< metal3 >>
rect 474 4216 1094 4221
rect 474 3916 484 4216
rect 1084 3916 1094 4216
rect 474 3911 1094 3916
rect 24106 4216 24726 4221
rect 24106 3916 24116 4216
rect 24716 3916 24726 4216
rect 24106 3911 24726 3916
rect 3998 3834 20878 3866
rect 3998 3620 4061 3834
rect 20846 3620 20878 3834
rect 3998 3600 20878 3620
rect 3998 3598 8352 3600
rect -15168 2940 -128 3086
rect -15168 2930 -974 2940
rect -15168 2240 -15016 2930
rect -14320 2242 -974 2930
rect -284 2242 -128 2940
rect -14320 2240 -128 2242
rect -15168 -10378 -128 2240
rect -15168 -10670 -13630 -10378
rect -2868 -10670 -128 -10378
rect -15168 -10978 -128 -10670
rect 2315 -10944 2413 -10939
rect 2314 -10945 2414 -10944
rect -15168 -11472 -1378 -10978
rect 2314 -11043 2315 -10945
rect 2413 -11043 2414 -10945
rect 2314 -11044 2414 -11043
rect 2315 -11049 2413 -11044
rect -15168 -11916 -1376 -11472
rect -1714 -11918 -1376 -11916
rect -8118 -26476 23968 -26430
rect -8118 -26630 -8072 -26476
rect 23928 -26630 23968 -26476
rect -8118 -26676 23968 -26630
rect -12226 -26816 -11606 -26811
rect -12226 -27116 -12216 -26816
rect -11616 -27116 -11606 -26816
rect -12226 -27121 -11606 -27116
rect 24206 -26816 24826 -26811
rect 24206 -27116 24216 -26816
rect 24816 -27116 24826 -26816
rect 24206 -27121 24826 -27116
<< via3 >>
rect 484 3916 1084 4216
rect 24116 3916 24716 4216
rect 4061 3620 20846 3834
rect -15016 2240 -14320 2930
rect -974 2242 -284 2940
rect 2315 -10949 2413 -10945
rect 2315 -11039 2319 -10949
rect 2319 -11039 2409 -10949
rect 2409 -11039 2413 -10949
rect 2315 -11043 2413 -11039
rect -8072 -26630 23928 -26476
rect -12216 -27116 -11616 -26816
rect 24216 -27116 24816 -26816
<< mimcap >>
rect -13982 2936 -7782 2986
rect -13982 2636 -8132 2936
rect -7832 2636 -7782 2936
rect -13982 2586 -7782 2636
rect -7582 2936 -1382 2986
rect -7582 2636 -1732 2936
rect -1432 2636 -1382 2936
rect -7582 2586 -1382 2636
rect -15068 1854 -14268 1904
rect -15068 -3846 -14618 1854
rect -14318 -3846 -14268 1854
rect -1024 1854 -224 1904
rect -13128 936 -7928 986
rect -13128 -3764 -8278 936
rect -7978 -3764 -7928 936
rect -13128 -3814 -7928 -3764
rect -7528 936 -2328 986
rect -7528 -3764 -2678 936
rect -2378 -3764 -2328 936
rect -7528 -3814 -2328 -3764
rect -15068 -3896 -14268 -3846
rect -1024 -3846 -574 1854
rect -274 -3846 -224 1854
rect -1024 -3896 -224 -3846
rect -15068 -4638 -14268 -4588
rect -15068 -10338 -14618 -4638
rect -14318 -10338 -14268 -4638
rect -13128 -4664 -7928 -4614
rect -13128 -9364 -8278 -4664
rect -7978 -9364 -7928 -4664
rect -13128 -9414 -7928 -9364
rect -7528 -4664 -2328 -4614
rect -7528 -9364 -2678 -4664
rect -2378 -9364 -2328 -4664
rect -7528 -9414 -2328 -9364
rect -1024 -4638 -224 -4588
rect -15068 -10388 -14268 -10338
rect -1024 -10338 -574 -4638
rect -274 -10338 -224 -4638
rect -1024 -10388 -224 -10338
rect -14482 -11064 -8282 -11014
rect -14482 -11364 -8632 -11064
rect -8332 -11364 -8282 -11064
rect -14482 -11414 -8282 -11364
rect -8082 -11064 -1882 -11014
rect -8082 -11364 -2232 -11064
rect -1932 -11364 -1882 -11064
rect -8082 -11414 -1882 -11364
<< mimcapcontact >>
rect -8132 2636 -7832 2936
rect -1732 2636 -1432 2936
rect -14618 -3846 -14318 1854
rect -8278 -3764 -7978 936
rect -2678 -3764 -2378 936
rect -574 -3846 -274 1854
rect -14618 -10338 -14318 -4638
rect -8278 -9364 -7978 -4664
rect -2678 -9364 -2378 -4664
rect -574 -10338 -274 -4638
rect -8632 -11364 -8332 -11064
rect -2232 -11364 -1932 -11064
<< metal4 >>
rect -15168 4216 25000 4400
rect -15168 3916 484 4216
rect 1084 3916 24116 4216
rect 24716 3916 25000 4216
rect -15168 3834 25000 3916
rect -15168 3620 4061 3834
rect 20846 3620 25000 3834
rect -15168 3600 25000 3620
rect -15168 2940 -128 3086
rect -15168 2936 -974 2940
rect -15168 2930 -8132 2936
rect -15168 2240 -15016 2930
rect -14320 2636 -8132 2930
rect -7832 2636 -1732 2936
rect -1432 2636 -974 2936
rect -14320 2242 -974 2636
rect -284 2242 -128 2940
rect -14320 2240 -128 2242
rect -15168 1910 -128 2240
rect -15168 1854 -13986 1910
rect -15168 -3846 -14618 1854
rect -14318 -3846 -13986 1854
rect -1428 1854 -128 1910
rect -15168 -4638 -13986 -3846
rect -15168 -10338 -14618 -4638
rect -14318 -10338 -13986 -4638
rect -13228 936 -2228 1086
rect -13228 -3764 -8278 936
rect -7978 -3764 -2678 936
rect -2378 -3764 -2228 936
rect -13228 -4664 -2228 -3764
rect -13228 -9364 -8278 -4664
rect -7978 -9364 -2678 -4664
rect -2378 -9364 -2228 -4664
rect -13228 -9816 -2228 -9364
rect -1428 -3846 -574 1854
rect -274 -3846 -128 1854
rect -1428 -4638 -128 -3846
rect -1428 -9436 -574 -4638
rect -13228 -9913 -1327 -9816
rect -13228 -9914 -2228 -9913
rect -15168 -10752 -13986 -10338
rect -15168 -10838 -2722 -10752
rect -15166 -10978 -2722 -10838
rect -15166 -11064 -1722 -10978
rect -15166 -11364 -8632 -11064
rect -8332 -11364 -2232 -11064
rect -1932 -11364 -1722 -11064
rect -15166 -11916 -1722 -11364
rect -1424 -11400 -1327 -9913
rect -1058 -10338 -574 -9436
rect -274 -10338 -128 -4638
rect -1058 -10848 -128 -10338
rect 226 -10945 2414 -10944
rect 226 -11043 2315 -10945
rect 2413 -11043 2414 -10945
rect 226 -11044 2414 -11043
rect 226 -11400 326 -11044
rect -1424 -11500 326 -11400
rect -15168 -26476 25000 -26400
rect -15168 -26630 -8072 -26476
rect 23928 -26630 25000 -26476
rect -15168 -26816 25000 -26630
rect -15168 -27116 -12216 -26816
rect -11616 -27116 24216 -26816
rect 24816 -27116 25000 -26816
rect -15168 -27200 25000 -27116
<< via4 >>
rect -15016 2240 -14320 2930
rect -974 2242 -284 2940
<< mimcap2 >>
rect -13982 2536 -8182 2986
rect -13982 2236 -13932 2536
rect -8232 2236 -8182 2536
rect -13982 2186 -8182 2236
rect -7582 2536 -1782 2986
rect -7582 2236 -7532 2536
rect -1832 2236 -1782 2536
rect -7582 2186 -1782 2236
rect -15068 -3946 -14668 1904
rect -15068 -4246 -15018 -3946
rect -14718 -4246 -14668 -3946
rect -13128 -3864 -8328 986
rect -13128 -4164 -13078 -3864
rect -8378 -4164 -8328 -3864
rect -13128 -4214 -8328 -4164
rect -7528 -3864 -2728 986
rect -7528 -4164 -7478 -3864
rect -2778 -4164 -2728 -3864
rect -7528 -4214 -2728 -4164
rect -1024 -3946 -624 1904
rect -15068 -4296 -14668 -4246
rect -1024 -4246 -974 -3946
rect -674 -4246 -624 -3946
rect -1024 -4296 -624 -4246
rect -15068 -10438 -14668 -4588
rect -13128 -9464 -8328 -4614
rect -13128 -9764 -13078 -9464
rect -8378 -9764 -8328 -9464
rect -13128 -9814 -8328 -9764
rect -7528 -9464 -2728 -4614
rect -7528 -9764 -7478 -9464
rect -2778 -9764 -2728 -9464
rect -7528 -9814 -2728 -9764
rect -15068 -10738 -15018 -10438
rect -14718 -10738 -14668 -10438
rect -15068 -10788 -14668 -10738
rect -1024 -10438 -624 -4588
rect -1024 -10724 -974 -10438
rect -674 -10724 -624 -10438
rect -1024 -10788 -624 -10724
rect -14482 -11464 -8682 -11014
rect -14482 -11764 -14432 -11464
rect -8732 -11764 -8682 -11464
rect -14482 -11814 -8682 -11764
rect -8082 -11464 -2282 -11014
rect -8082 -11764 -8032 -11464
rect -2332 -11764 -2282 -11464
rect -8082 -11814 -2282 -11764
<< mimcap2contact >>
rect -13932 2236 -8232 2536
rect -7532 2236 -1832 2536
rect -15018 -4246 -14718 -3946
rect -13078 -4164 -8378 -3864
rect -7478 -4164 -2778 -3864
rect -974 -4246 -674 -3946
rect -13078 -9764 -8378 -9464
rect -7478 -9764 -2778 -9464
rect -15018 -10738 -14718 -10438
rect -974 -10724 -674 -10438
rect -14432 -11764 -8732 -11464
rect -8032 -11764 -2332 -11464
<< metal5 >>
rect -15168 2940 -128 3086
rect -15168 2930 -974 2940
rect -15168 2240 -15016 2930
rect -14320 2536 -974 2930
rect -14320 2240 -13932 2536
rect -15168 2236 -13932 2240
rect -8232 2236 -7532 2536
rect -1832 2242 -974 2536
rect -284 2242 -128 2940
rect -1832 2236 -128 2242
rect -15168 -3864 -128 2236
rect -15168 -3946 -13078 -3864
rect -15168 -4246 -15018 -3946
rect -14718 -4164 -13078 -3946
rect -8378 -4164 -7478 -3864
rect -2778 -3946 -128 -3864
rect -2778 -4164 -974 -3946
rect -14718 -4246 -974 -4164
rect -674 -4246 -128 -3946
rect -15168 -9464 -128 -4246
rect -15168 -9764 -13078 -9464
rect -8378 -9764 -7478 -9464
rect -2778 -9764 -128 -9464
rect -15168 -10438 -128 -9764
rect -15168 -10738 -15018 -10438
rect -14718 -10724 -974 -10438
rect -674 -10724 -128 -10438
rect -14718 -10738 -128 -10724
rect -15168 -10764 -128 -10738
rect -15168 -11464 -130 -10764
rect -15168 -11764 -14432 -11464
rect -8732 -11764 -8032 -11464
rect -2332 -11764 -130 -11464
rect -15168 -11916 -130 -11764
use ptap  ptap_251 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/ptap
timestamp 1624298412
transform 1 0 -10304 0 1 -26298
box 70 126 186 240
use ptap  ptap_253
timestamp 1624298412
transform 1 0 -9286 0 1 -26298
box 70 126 186 240
use ptap  ptap_252
timestamp 1624298412
transform 1 0 -8268 0 1 -26298
box 70 126 186 240
use ptap  ptap_255
timestamp 1624298412
transform 1 0 -7250 0 1 -26298
box 70 126 186 240
use ptap  ptap_254
timestamp 1624298412
transform 1 0 -6232 0 1 -26298
box 70 126 186 240
use ptap  ptap_257
timestamp 1624298412
transform 1 0 -5214 0 1 -26298
box 70 126 186 240
use ptap  ptap_256
timestamp 1624298412
transform 1 0 -4196 0 1 -26298
box 70 126 186 240
use ptap  ptap_259
timestamp 1624298412
transform 1 0 -3178 0 1 -26298
box 70 126 186 240
use ptap  ptap_258
timestamp 1624298412
transform 1 0 -2160 0 1 -26298
box 70 126 186 240
use ptap  ptap_261
timestamp 1624298412
transform 1 0 -1142 0 1 -26298
box 70 126 186 240
use ptap  ptap_260
timestamp 1624298412
transform 1 0 -124 0 1 -26298
box 70 126 186 240
use ptap  ptap_234
timestamp 1624298412
transform 1 0 2986 0 1 -26380
box 70 126 186 240
use ptap  ptap_235
timestamp 1624298412
transform 1 0 4004 0 1 -26380
box 70 126 186 240
use ptap  ptap_236
timestamp 1624298412
transform 1 0 5022 0 1 -26380
box 70 126 186 240
use ptap  ptap_237
timestamp 1624298412
transform 1 0 6040 0 1 -26380
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_FYXD5N  sky130_fd_pr__nfet_01v8_FYXD5N_0
timestamp 1624298412
transform 1 0 -4943 0 1 -25440
box -5119 -388 5119 388
use ptap  ptap_238
timestamp 1624298412
transform 1 0 7058 0 1 -26380
box 70 126 186 240
use ptap  ptap_239
timestamp 1624298412
transform 1 0 8076 0 1 -26380
box 70 126 186 240
use ptap  ptap_220
timestamp 1624298412
transform 1 0 9094 0 1 -26380
box 70 126 186 240
use ptap  ptap_221
timestamp 1624298412
transform 1 0 10112 0 1 -26380
box 70 126 186 240
use ptap  ptap_222
timestamp 1624298412
transform 1 0 11130 0 1 -26380
box 70 126 186 240
use ptap  ptap_223
timestamp 1624298412
transform 1 0 12148 0 1 -26380
box 70 126 186 240
use ptap  ptap_224
timestamp 1624298412
transform 1 0 13166 0 1 -26380
box 70 126 186 240
use ptap  ptap_225
timestamp 1624298412
transform 1 0 14184 0 1 -26380
box 70 126 186 240
use ptap  ptap_226
timestamp 1624298412
transform 1 0 15202 0 1 -26380
box 70 126 186 240
use ptap  ptap_227
timestamp 1624298412
transform 1 0 16220 0 1 -26380
box 70 126 186 240
use ptap  ptap_228
timestamp 1624298412
transform 1 0 17238 0 1 -26380
box 70 126 186 240
use ptap  ptap_229
timestamp 1624298412
transform 1 0 18256 0 1 -26380
box 70 126 186 240
use ptap  ptap_230
timestamp 1624298412
transform 1 0 19274 0 1 -26380
box 70 126 186 240
use ptap  ptap_231
timestamp 1624298412
transform 1 0 20292 0 1 -26380
box 70 126 186 240
use ptap  ptap_232
timestamp 1624298412
transform 1 0 21310 0 1 -26380
box 70 126 186 240
use ptap  ptap_233
timestamp 1624298412
transform 1 0 22328 0 1 -26380
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_6
timestamp 1624298412
transform -1 0 12777 0 -1 -25630
box -10209 -388 10209 388
use ptap  ptap_240
timestamp 1624298412
transform 1 0 -10114 0 1 -24852
box 70 126 186 240
use ptap  ptap_242
timestamp 1624298412
transform 1 0 -9096 0 1 -24852
box 70 126 186 240
use ptap  ptap_241
timestamp 1624298412
transform 1 0 -8078 0 1 -24852
box 70 126 186 240
use ptap  ptap_244
timestamp 1624298412
transform 1 0 -7060 0 1 -24852
box 70 126 186 240
use ptap  ptap_243
timestamp 1624298412
transform 1 0 -6042 0 1 -24852
box 70 126 186 240
use ptap  ptap_246
timestamp 1624298412
transform 1 0 -5024 0 1 -24852
box 70 126 186 240
use ptap  ptap_245
timestamp 1624298412
transform 1 0 -4006 0 1 -24852
box 70 126 186 240
use ptap  ptap_247
timestamp 1624298412
transform 1 0 -1970 0 1 -24852
box 70 126 186 240
use ptap  ptap_248
timestamp 1624298412
transform 1 0 -2988 0 1 -24852
box 70 126 186 240
use ptap  ptap_250
timestamp 1624298412
transform 1 0 -952 0 1 -24852
box 70 126 186 240
use ptap  ptap_249
timestamp 1624298412
transform 1 0 66 0 1 -24852
box 70 126 186 240
use ptap  ptap_214
timestamp 1624298412
transform 1 0 2998 0 1 -25202
box 70 126 186 240
use ptap  ptap_215
timestamp 1624298412
transform 1 0 4016 0 1 -25202
box 70 126 186 240
use ptap  ptap_216
timestamp 1624298412
transform 1 0 5034 0 1 -25202
box 70 126 186 240
use ptap  ptap_217
timestamp 1624298412
transform 1 0 6052 0 1 -25202
box 70 126 186 240
use ptap  ptap_218
timestamp 1624298412
transform 1 0 7070 0 1 -25202
box 70 126 186 240
use ptap  ptap_219
timestamp 1624298412
transform 1 0 8088 0 1 -25202
box 70 126 186 240
use ptap  ptap_200
timestamp 1624298412
transform 1 0 9106 0 1 -25202
box 70 126 186 240
use ptap  ptap_201
timestamp 1624298412
transform 1 0 10124 0 1 -25202
box 70 126 186 240
use ptap  ptap_202
timestamp 1624298412
transform 1 0 11142 0 1 -25202
box 70 126 186 240
use ptap  ptap_204
timestamp 1624298412
transform 1 0 13178 0 1 -25202
box 70 126 186 240
use ptap  ptap_203
timestamp 1624298412
transform 1 0 12160 0 1 -25202
box 70 126 186 240
use ptap  ptap_205
timestamp 1624298412
transform 1 0 14196 0 1 -25202
box 70 126 186 240
use ptap  ptap_206
timestamp 1624298412
transform 1 0 15214 0 1 -25202
box 70 126 186 240
use ptap  ptap_207
timestamp 1624298412
transform 1 0 16232 0 1 -25202
box 70 126 186 240
use ptap  ptap_208
timestamp 1624298412
transform 1 0 17250 0 1 -25202
box 70 126 186 240
use ptap  ptap_209
timestamp 1624298412
transform 1 0 18268 0 1 -25202
box 70 126 186 240
use ptap  ptap_210
timestamp 1624298412
transform 1 0 19286 0 1 -25202
box 70 126 186 240
use ptap  ptap_211
timestamp 1624298412
transform 1 0 20304 0 1 -25202
box 70 126 186 240
use ptap  ptap_212
timestamp 1624298412
transform 1 0 21322 0 1 -25202
box 70 126 186 240
use ptap  ptap_213
timestamp 1624298412
transform 1 0 22340 0 1 -25202
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_9
timestamp 1624298412
transform 1 0 12777 0 1 -24398
box -10209 -388 10209 388
use sky130_fd_pr__nfet_01v8_lvt_ZYX5GY  sky130_fd_pr__nfet_01v8_lvt_ZYX5GY_3
timestamp 1624298412
transform 1 0 -4892 0 1 -23898
box -5628 -388 5628 388
use ptap  ptap_197
timestamp 1624298412
transform 1 0 6040 0 1 -23956
box 70 126 186 240
use ptap  ptap_196
timestamp 1624298412
transform 1 0 5022 0 1 -23956
box 70 126 186 240
use ptap  ptap_195
timestamp 1624298412
transform 1 0 4004 0 1 -23956
box 70 126 186 240
use ptap  ptap_194
timestamp 1624298412
transform 1 0 2986 0 1 -23956
box 70 126 186 240
use ptap  ptap_264
timestamp 1624298412
transform 1 0 -9096 0 1 -23510
box 70 126 186 240
use ptap  ptap_262
timestamp 1624298412
transform 1 0 -10114 0 1 -23510
box 70 126 186 240
use ptap  ptap_263
timestamp 1624298412
transform 1 0 -8078 0 1 -23510
box 70 126 186 240
use ptap  ptap_266
timestamp 1624298412
transform 1 0 -7060 0 1 -23510
box 70 126 186 240
use ptap  ptap_265
timestamp 1624298412
transform 1 0 -6042 0 1 -23510
box 70 126 186 240
use ptap  ptap_268
timestamp 1624298412
transform 1 0 -5024 0 1 -23510
box 70 126 186 240
use ptap  ptap_270
timestamp 1624298412
transform 1 0 -2988 0 1 -23510
box 70 126 186 240
use ptap  ptap_267
timestamp 1624298412
transform 1 0 -4006 0 1 -23510
box 70 126 186 240
use ptap  ptap_269
timestamp 1624298412
transform 1 0 -1970 0 1 -23510
box 70 126 186 240
use ptap  ptap_272
timestamp 1624298412
transform 1 0 -952 0 1 -23510
box 70 126 186 240
use ptap  ptap_271
timestamp 1624298412
transform 1 0 66 0 1 -23510
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_lvt_ZYX5GY  sky130_fd_pr__nfet_01v8_lvt_ZYX5GY_2
timestamp 1624298412
transform 1 0 -4892 0 1 -22786
box -5628 -388 5628 388
use ptap  ptap_198
timestamp 1624298412
transform 1 0 7058 0 1 -23956
box 70 126 186 240
use ptap  ptap_199
timestamp 1624298412
transform 1 0 8076 0 1 -23956
box 70 126 186 240
use ptap  ptap_180
timestamp 1624298412
transform 1 0 9094 0 1 -23956
box 70 126 186 240
use ptap  ptap_181
timestamp 1624298412
transform 1 0 10112 0 1 -23956
box 70 126 186 240
use ptap  ptap_182
timestamp 1624298412
transform 1 0 11130 0 1 -23956
box 70 126 186 240
use ptap  ptap_183
timestamp 1624298412
transform 1 0 12148 0 1 -23956
box 70 126 186 240
use ptap  ptap_184
timestamp 1624298412
transform 1 0 13166 0 1 -23956
box 70 126 186 240
use ptap  ptap_185
timestamp 1624298412
transform 1 0 14184 0 1 -23956
box 70 126 186 240
use ptap  ptap_186
timestamp 1624298412
transform 1 0 15202 0 1 -23956
box 70 126 186 240
use ptap  ptap_187
timestamp 1624298412
transform 1 0 16220 0 1 -23956
box 70 126 186 240
use ptap  ptap_188
timestamp 1624298412
transform 1 0 17238 0 1 -23956
box 70 126 186 240
use ptap  ptap_189
timestamp 1624298412
transform 1 0 18256 0 1 -23956
box 70 126 186 240
use ptap  ptap_190
timestamp 1624298412
transform 1 0 19274 0 1 -23956
box 70 126 186 240
use ptap  ptap_191
timestamp 1624298412
transform 1 0 20292 0 1 -23956
box 70 126 186 240
use ptap  ptap_192
timestamp 1624298412
transform 1 0 21310 0 1 -23956
box 70 126 186 240
use ptap  ptap_193
timestamp 1624298412
transform 1 0 22328 0 1 -23956
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_5
timestamp 1624298412
transform 1 0 12777 0 1 -23164
box -10209 -388 10209 388
use ptap  ptap_273
timestamp 1624298412
transform 1 0 -10114 0 1 -22404
box 70 126 186 240
use ptap  ptap_275
timestamp 1624298412
transform 1 0 -9096 0 1 -22404
box 70 126 186 240
use ptap  ptap_274
timestamp 1624298412
transform 1 0 -8078 0 1 -22404
box 70 126 186 240
use ptap  ptap_277
timestamp 1624298412
transform 1 0 -7060 0 1 -22404
box 70 126 186 240
use ptap  ptap_276
timestamp 1624298412
transform 1 0 -6042 0 1 -22404
box 70 126 186 240
use ptap  ptap_279
timestamp 1624298412
transform 1 0 -5024 0 1 -22404
box 70 126 186 240
use ptap  ptap_278
timestamp 1624298412
transform 1 0 -4006 0 1 -22404
box 70 126 186 240
use ptap  ptap_280
timestamp 1624298412
transform 1 0 -1970 0 1 -22404
box 70 126 186 240
use ptap  ptap_281
timestamp 1624298412
transform 1 0 -2988 0 1 -22404
box 70 126 186 240
use ptap  ptap_283
timestamp 1624298412
transform 1 0 -952 0 1 -22404
box 70 126 186 240
use ptap  ptap_282
timestamp 1624298412
transform 1 0 66 0 1 -22404
box 70 126 186 240
use ptap  ptap_174
timestamp 1624298412
transform 1 0 2986 0 1 -22720
box 70 126 186 240
use ptap  ptap_175
timestamp 1624298412
transform 1 0 4004 0 1 -22720
box 70 126 186 240
use ptap  ptap_176
timestamp 1624298412
transform 1 0 5022 0 1 -22720
box 70 126 186 240
use ptap  ptap_177
timestamp 1624298412
transform 1 0 6040 0 1 -22720
box 70 126 186 240
use ptap  ptap_178
timestamp 1624298412
transform 1 0 7058 0 1 -22720
box 70 126 186 240
use ptap  ptap_179
timestamp 1624298412
transform 1 0 8076 0 1 -22720
box 70 126 186 240
use ptap  ptap_160
timestamp 1624298412
transform 1 0 9094 0 1 -22720
box 70 126 186 240
use ptap  ptap_161
timestamp 1624298412
transform 1 0 10112 0 1 -22720
box 70 126 186 240
use ptap  ptap_162
timestamp 1624298412
transform 1 0 11130 0 1 -22720
box 70 126 186 240
use ptap  ptap_164
timestamp 1624298412
transform 1 0 13166 0 1 -22720
box 70 126 186 240
use ptap  ptap_163
timestamp 1624298412
transform 1 0 12148 0 1 -22720
box 70 126 186 240
use ptap  ptap_165
timestamp 1624298412
transform 1 0 14184 0 1 -22720
box 70 126 186 240
use ptap  ptap_166
timestamp 1624298412
transform 1 0 15202 0 1 -22720
box 70 126 186 240
use ptap  ptap_167
timestamp 1624298412
transform 1 0 16220 0 1 -22720
box 70 126 186 240
use ptap  ptap_168
timestamp 1624298412
transform 1 0 17238 0 1 -22720
box 70 126 186 240
use ptap  ptap_169
timestamp 1624298412
transform 1 0 18256 0 1 -22720
box 70 126 186 240
use ptap  ptap_170
timestamp 1624298412
transform 1 0 19274 0 1 -22720
box 70 126 186 240
use ptap  ptap_171
timestamp 1624298412
transform 1 0 20292 0 1 -22720
box 70 126 186 240
use ptap  ptap_172
timestamp 1624298412
transform 1 0 21310 0 1 -22720
box 70 126 186 240
use ptap  ptap_173
timestamp 1624298412
transform 1 0 22328 0 1 -22720
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_4
timestamp 1624298412
transform 1 0 12777 0 1 -21932
box -10209 -388 10209 388
use sky130_fd_pr__nfet_01v8_lvt_ZYX5GY  sky130_fd_pr__nfet_01v8_lvt_ZYX5GY_1
timestamp 1624298412
transform 1 0 -4892 0 1 -21674
box -5628 -388 5628 388
use ptap  ptap_284
timestamp 1624298412
transform 1 0 -10092 0 1 -21296
box 70 126 186 240
use ptap  ptap_286
timestamp 1624298412
transform 1 0 -9074 0 1 -21296
box 70 126 186 240
use ptap  ptap_285
timestamp 1624298412
transform 1 0 -8056 0 1 -21296
box 70 126 186 240
use ptap  ptap_288
timestamp 1624298412
transform 1 0 -7038 0 1 -21296
box 70 126 186 240
use ptap  ptap_287
timestamp 1624298412
transform 1 0 -6020 0 1 -21296
box 70 126 186 240
use ptap  ptap_290
timestamp 1624298412
transform 1 0 -5002 0 1 -21296
box 70 126 186 240
use ptap  ptap_289
timestamp 1624298412
transform 1 0 -3984 0 1 -21296
box 70 126 186 240
use ptap  ptap_292
timestamp 1624298412
transform 1 0 -2966 0 1 -21296
box 70 126 186 240
use ptap  ptap_291
timestamp 1624298412
transform 1 0 -1948 0 1 -21296
box 70 126 186 240
use ptap  ptap_294
timestamp 1624298412
transform 1 0 -930 0 1 -21296
box 70 126 186 240
use ptap  ptap_293
timestamp 1624298412
transform 1 0 88 0 1 -21296
box 70 126 186 240
use ptap  ptap_154
timestamp 1624298412
transform 1 0 2974 0 1 -21496
box 70 126 186 240
use ptap  ptap_155
timestamp 1624298412
transform 1 0 3992 0 1 -21496
box 70 126 186 240
use ptap  ptap_156
timestamp 1624298412
transform 1 0 5010 0 1 -21496
box 70 126 186 240
use ptap  ptap_157
timestamp 1624298412
transform 1 0 6028 0 1 -21496
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_lvt_ZYX5GY  sky130_fd_pr__nfet_01v8_lvt_ZYX5GY_0
timestamp 1624298412
transform 1 0 -4892 0 1 -20562
box -5628 -388 5628 388
use ptap  ptap_158
timestamp 1624298412
transform 1 0 7046 0 1 -21496
box 70 126 186 240
use ptap  ptap_159
timestamp 1624298412
transform 1 0 8064 0 1 -21496
box 70 126 186 240
use ptap  ptap_140
timestamp 1624298412
transform 1 0 9082 0 1 -21496
box 70 126 186 240
use ptap  ptap_141
timestamp 1624298412
transform 1 0 10100 0 1 -21496
box 70 126 186 240
use ptap  ptap_142
timestamp 1624298412
transform 1 0 11118 0 1 -21496
box 70 126 186 240
use ptap  ptap_143
timestamp 1624298412
transform 1 0 12136 0 1 -21496
box 70 126 186 240
use ptap  ptap_144
timestamp 1624298412
transform 1 0 13154 0 1 -21496
box 70 126 186 240
use ptap  ptap_145
timestamp 1624298412
transform 1 0 14172 0 1 -21496
box 70 126 186 240
use ptap  ptap_146
timestamp 1624298412
transform 1 0 15190 0 1 -21496
box 70 126 186 240
use ptap  ptap_147
timestamp 1624298412
transform 1 0 16208 0 1 -21496
box 70 126 186 240
use ptap  ptap_148
timestamp 1624298412
transform 1 0 17226 0 1 -21496
box 70 126 186 240
use ptap  ptap_149
timestamp 1624298412
transform 1 0 18244 0 1 -21496
box 70 126 186 240
use ptap  ptap_150
timestamp 1624298412
transform 1 0 19262 0 1 -21496
box 70 126 186 240
use ptap  ptap_151
timestamp 1624298412
transform 1 0 20280 0 1 -21496
box 70 126 186 240
use ptap  ptap_152
timestamp 1624298412
transform 1 0 21298 0 1 -21496
box 70 126 186 240
use ptap  ptap_153
timestamp 1624298412
transform 1 0 22316 0 1 -21496
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_3
timestamp 1624298412
transform 1 0 12777 0 1 -20698
box -10209 -388 10209 388
use ptap  ptap_295
timestamp 1624298412
transform 1 0 -10104 0 1 -20154
box 70 126 186 240
use ptap  ptap_297
timestamp 1624298412
transform 1 0 -9086 0 1 -20154
box 70 126 186 240
use ptap  ptap_296
timestamp 1624298412
transform 1 0 -8068 0 1 -20154
box 70 126 186 240
use ptap  ptap_299
timestamp 1624298412
transform 1 0 -7050 0 1 -20154
box 70 126 186 240
use ptap  ptap_298
timestamp 1624298412
transform 1 0 -6032 0 1 -20154
box 70 126 186 240
use ptap  ptap_301
timestamp 1624298412
transform 1 0 -5014 0 1 -20154
box 70 126 186 240
use ptap  ptap_300
timestamp 1624298412
transform 1 0 -3996 0 1 -20154
box 70 126 186 240
use ptap  ptap_303
timestamp 1624298412
transform 1 0 -2978 0 1 -20154
box 70 126 186 240
use ptap  ptap_302
timestamp 1624298412
transform 1 0 -1960 0 1 -20154
box 70 126 186 240
use ptap  ptap_305
timestamp 1624298412
transform 1 0 -942 0 1 -20154
box 70 126 186 240
use ptap  ptap_304
timestamp 1624298412
transform 1 0 76 0 1 -20154
box 70 126 186 240
use ptap  ptap_134
timestamp 1624298412
transform 1 0 2998 0 1 -20260
box 70 126 186 240
use ptap  ptap_135
timestamp 1624298412
transform 1 0 4016 0 1 -20260
box 70 126 186 240
use ptap  ptap_136
timestamp 1624298412
transform 1 0 5034 0 1 -20260
box 70 126 186 240
use ptap  ptap_137
timestamp 1624298412
transform 1 0 6052 0 1 -20260
box 70 126 186 240
use ptap  ptap_138
timestamp 1624298412
transform 1 0 7070 0 1 -20260
box 70 126 186 240
use ptap  ptap_139
timestamp 1624298412
transform 1 0 8088 0 1 -20260
box 70 126 186 240
use ptap  ptap_120
timestamp 1624298412
transform 1 0 9106 0 1 -20260
box 70 126 186 240
use ptap  ptap_121
timestamp 1624298412
transform 1 0 10124 0 1 -20260
box 70 126 186 240
use ptap  ptap_122
timestamp 1624298412
transform 1 0 11142 0 1 -20260
box 70 126 186 240
use ptap  ptap_123
timestamp 1624298412
transform 1 0 12160 0 1 -20260
box 70 126 186 240
use ptap  ptap_124
timestamp 1624298412
transform 1 0 13178 0 1 -20260
box 70 126 186 240
use ptap  ptap_125
timestamp 1624298412
transform 1 0 14196 0 1 -20260
box 70 126 186 240
use ptap  ptap_126
timestamp 1624298412
transform 1 0 15214 0 1 -20260
box 70 126 186 240
use ptap  ptap_127
timestamp 1624298412
transform 1 0 16232 0 1 -20260
box 70 126 186 240
use ptap  ptap_128
timestamp 1624298412
transform 1 0 17250 0 1 -20260
box 70 126 186 240
use ptap  ptap_129
timestamp 1624298412
transform 1 0 18268 0 1 -20260
box 70 126 186 240
use ptap  ptap_130
timestamp 1624298412
transform 1 0 19286 0 1 -20260
box 70 126 186 240
use ptap  ptap_131
timestamp 1624298412
transform 1 0 20304 0 1 -20260
box 70 126 186 240
use ptap  ptap_132
timestamp 1624298412
transform 1 0 21322 0 1 -20260
box 70 126 186 240
use ptap  ptap_133
timestamp 1624298412
transform 1 0 22340 0 1 -20260
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_2
timestamp 1624298412
transform 1 0 12777 0 1 -19464
box -10209 -388 10209 388
use ptap  ptap_318
timestamp 1624298412
transform 1 0 -8290 0 1 -19206
box 70 126 186 240
use ptap  ptap_317
timestamp 1624298412
transform 1 0 -7272 0 1 -19206
box 70 126 186 240
use ptap  ptap_316
timestamp 1624298412
transform 1 0 -9308 0 1 -19206
box 70 126 186 240
use ptap  ptap_319
timestamp 1624298412
transform 1 0 -5236 0 1 -19206
box 70 126 186 240
use ptap  ptap_320
timestamp 1624298412
transform 1 0 -6254 0 1 -19206
box 70 126 186 240
use ptap  ptap_322
timestamp 1624298412
transform 1 0 -4218 0 1 -19206
box 70 126 186 240
use ptap  ptap_321
timestamp 1624298412
transform 1 0 -3200 0 1 -19206
box 70 126 186 240
use ptap  ptap_323
timestamp 1624298412
transform 1 0 -1164 0 1 -19206
box 70 126 186 240
use ptap  ptap_324
timestamp 1624298412
transform 1 0 -2182 0 1 -19206
box 70 126 186 240
use ptap  ptap_325
timestamp 1624298412
transform 1 0 -136 0 1 -19206
box 70 126 186 240
use ptap  ptap_114
timestamp 1624298412
transform 1 0 2998 0 1 -19012
box 70 126 186 240
use ptap  ptap_115
timestamp 1624298412
transform 1 0 4016 0 1 -19012
box 70 126 186 240
use ptap  ptap_116
timestamp 1624298412
transform 1 0 5034 0 1 -19012
box 70 126 186 240
use ptap  ptap_117
timestamp 1624298412
transform 1 0 6052 0 1 -19012
box 70 126 186 240
use ptap  ptap_118
timestamp 1624298412
transform 1 0 7070 0 1 -19012
box 70 126 186 240
use ptap  ptap_100
timestamp 1624298412
transform 1 0 9106 0 1 -19012
box 70 126 186 240
use ptap  ptap_119
timestamp 1624298412
transform 1 0 8088 0 1 -19012
box 70 126 186 240
use ptap  ptap_101
timestamp 1624298412
transform 1 0 10124 0 1 -19012
box 70 126 186 240
use ptap  ptap_102
timestamp 1624298412
transform 1 0 11142 0 1 -19012
box 70 126 186 240
use ptap  ptap_103
timestamp 1624298412
transform 1 0 12160 0 1 -19012
box 70 126 186 240
use ptap  ptap_104
timestamp 1624298412
transform 1 0 13178 0 1 -19012
box 70 126 186 240
use ptap  ptap_105
timestamp 1624298412
transform 1 0 14196 0 1 -19012
box 70 126 186 240
use ptap  ptap_106
timestamp 1624298412
transform 1 0 15214 0 1 -19012
box 70 126 186 240
use ptap  ptap_107
timestamp 1624298412
transform 1 0 16232 0 1 -19012
box 70 126 186 240
use ptap  ptap_108
timestamp 1624298412
transform 1 0 17250 0 1 -19012
box 70 126 186 240
use ptap  ptap_109
timestamp 1624298412
transform 1 0 18268 0 1 -19012
box 70 126 186 240
use ptap  ptap_110
timestamp 1624298412
transform 1 0 19286 0 1 -19012
box 70 126 186 240
use ptap  ptap_111
timestamp 1624298412
transform 1 0 20304 0 1 -19012
box 70 126 186 240
use ptap  ptap_112
timestamp 1624298412
transform 1 0 21322 0 1 -19012
box 70 126 186 240
use ptap  ptap_113
timestamp 1624298412
transform 1 0 22340 0 1 -19012
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_1
timestamp 1624298412
transform 1 0 12777 0 1 -18232
box -10209 -388 10209 388
use ptap  ptap_314
timestamp 1624298412
transform 1 0 -8278 0 1 -18312
box 70 126 186 240
use ptap  ptap_313
timestamp 1624298412
transform 1 0 -7260 0 1 -18312
box 70 126 186 240
use ptap  ptap_315
timestamp 1624298412
transform 1 0 -9296 0 1 -18312
box 70 126 186 240
use ptap  ptap_310
timestamp 1624298412
transform 1 0 -4206 0 1 -18312
box 70 126 186 240
use ptap  ptap_311
timestamp 1624298412
transform 1 0 -5224 0 1 -18312
box 70 126 186 240
use ptap  ptap_312
timestamp 1624298412
transform 1 0 -6242 0 1 -18312
box 70 126 186 240
use ptap  ptap_307
timestamp 1624298412
transform 1 0 -1152 0 1 -18312
box 70 126 186 240
use ptap  ptap_308
timestamp 1624298412
transform 1 0 -2170 0 1 -18312
box 70 126 186 240
use ptap  ptap_309
timestamp 1624298412
transform 1 0 -3188 0 1 -18312
box 70 126 186 240
use ptap  ptap_306
timestamp 1624298412
transform 1 0 -124 0 1 -18312
box 70 126 186 240
use ptap  ptap_94
timestamp 1624298412
transform 1 0 2986 0 1 -17776
box 70 126 186 240
use ptap  ptap_95
timestamp 1624298412
transform 1 0 4004 0 1 -17776
box 70 126 186 240
use ptap  ptap_96
timestamp 1624298412
transform 1 0 5022 0 1 -17776
box 70 126 186 240
use ptap  ptap_97
timestamp 1624298412
transform 1 0 6040 0 1 -17776
box 70 126 186 240
use ptap  ptap_98
timestamp 1624298412
transform 1 0 7058 0 1 -17776
box 70 126 186 240
use ptap  ptap_80
timestamp 1624298412
transform 1 0 9094 0 1 -17776
box 70 126 186 240
use ptap  ptap_99
timestamp 1624298412
transform 1 0 8076 0 1 -17776
box 70 126 186 240
use ptap  ptap_81
timestamp 1624298412
transform 1 0 10112 0 1 -17776
box 70 126 186 240
use ptap  ptap_82
timestamp 1624298412
transform 1 0 11130 0 1 -17776
box 70 126 186 240
use ptap  ptap_83
timestamp 1624298412
transform 1 0 12148 0 1 -17776
box 70 126 186 240
use ptap  ptap_85
timestamp 1624298412
transform 1 0 14184 0 1 -17776
box 70 126 186 240
use ptap  ptap_84
timestamp 1624298412
transform 1 0 13166 0 1 -17776
box 70 126 186 240
use ptap  ptap_86
timestamp 1624298412
transform 1 0 15202 0 1 -17776
box 70 126 186 240
use ptap  ptap_87
timestamp 1624298412
transform 1 0 16220 0 1 -17776
box 70 126 186 240
use ptap  ptap_88
timestamp 1624298412
transform 1 0 17238 0 1 -17776
box 70 126 186 240
use ptap  ptap_90
timestamp 1624298412
transform 1 0 19274 0 1 -17776
box 70 126 186 240
use ptap  ptap_89
timestamp 1624298412
transform 1 0 18256 0 1 -17776
box 70 126 186 240
use ptap  ptap_91
timestamp 1624298412
transform 1 0 20292 0 1 -17776
box 70 126 186 240
use ptap  ptap_92
timestamp 1624298412
transform 1 0 21310 0 1 -17776
box 70 126 186 240
use ptap  ptap_93
timestamp 1624298412
transform 1 0 22328 0 1 -17776
box 70 126 186 240
use ptap  ptap_326
timestamp 1624298412
transform 1 0 -9296 0 1 -17494
box 70 126 186 240
use ptap  ptap_328
timestamp 1624298412
transform 1 0 -7260 0 1 -17494
box 70 126 186 240
use ptap  ptap_327
timestamp 1624298412
transform 1 0 -8278 0 1 -17494
box 70 126 186 240
use ptap  ptap_330
timestamp 1624298412
transform 1 0 -5224 0 1 -17494
box 70 126 186 240
use ptap  ptap_329
timestamp 1624298412
transform 1 0 -6242 0 1 -17494
box 70 126 186 240
use ptap  ptap_331
timestamp 1624298412
transform 1 0 -4206 0 1 -17494
box 70 126 186 240
use ptap  ptap_333
timestamp 1624298412
transform 1 0 -2170 0 1 -17494
box 70 126 186 240
use ptap  ptap_332
timestamp 1624298412
transform 1 0 -3188 0 1 -17494
box 70 126 186 240
use ptap  ptap_334
timestamp 1624298412
transform 1 0 -1152 0 1 -17494
box 70 126 186 240
use ptap  ptap_335
timestamp 1624298412
transform 1 0 -124 0 1 -17494
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_0
timestamp 1624298412
transform 1 0 12777 0 1 -16998
box -10209 -388 10209 388
use sky130_fd_pr__nfet_01v8_lvt_XH9Q8F  sky130_fd_pr__nfet_01v8_lvt_XH9Q8F_1
timestamp 1624298412
transform 1 0 -4586 0 1 -17311
box -4610 -1615 4610 1615
use ptap  ptap_336
timestamp 1624298412
transform 1 0 -9296 0 1 -16676
box 70 126 186 240
use ptap  ptap_338
timestamp 1624298412
transform 1 0 -7260 0 1 -16676
box 70 126 186 240
use ptap  ptap_337
timestamp 1624298412
transform 1 0 -8278 0 1 -16676
box 70 126 186 240
use ptap  ptap_339
timestamp 1624298412
transform 1 0 -6242 0 1 -16676
box 70 126 186 240
use ptap  ptap_340
timestamp 1624298412
transform 1 0 -5224 0 1 -16676
box 70 126 186 240
use ptap  ptap_341
timestamp 1624298412
transform 1 0 -4206 0 1 -16676
box 70 126 186 240
use ptap  ptap_342
timestamp 1624298412
transform 1 0 -3188 0 1 -16676
box 70 126 186 240
use ptap  ptap_343
timestamp 1624298412
transform 1 0 -2170 0 1 -16676
box 70 126 186 240
use ptap  ptap_344
timestamp 1624298412
transform 1 0 -1152 0 1 -16676
box 70 126 186 240
use ptap  ptap_345
timestamp 1624298412
transform 1 0 -124 0 1 -16676
box 70 126 186 240
use ptap  ptap_74
timestamp 1624298412
transform 1 0 2986 0 1 -16552
box 70 126 186 240
use ptap  ptap_75
timestamp 1624298412
transform 1 0 4004 0 1 -16552
box 70 126 186 240
use ptap  ptap_76
timestamp 1624298412
transform 1 0 5022 0 1 -16552
box 70 126 186 240
use ptap  ptap_77
timestamp 1624298412
transform 1 0 6040 0 1 -16552
box 70 126 186 240
use ptap  ptap_78
timestamp 1624298412
transform 1 0 7058 0 1 -16552
box 70 126 186 240
use ptap  ptap_79
timestamp 1624298412
transform 1 0 8076 0 1 -16552
box 70 126 186 240
use ptap  ptap_60
timestamp 1624298412
transform 1 0 9094 0 1 -16552
box 70 126 186 240
use ptap  ptap_61
timestamp 1624298412
transform 1 0 10112 0 1 -16552
box 70 126 186 240
use ptap  ptap_62
timestamp 1624298412
transform 1 0 11130 0 1 -16552
box 70 126 186 240
use ptap  ptap_63
timestamp 1624298412
transform 1 0 12148 0 1 -16552
box 70 126 186 240
use ptap  ptap_64
timestamp 1624298412
transform 1 0 13166 0 1 -16552
box 70 126 186 240
use ptap  ptap_65
timestamp 1624298412
transform 1 0 14184 0 1 -16552
box 70 126 186 240
use ptap  ptap_66
timestamp 1624298412
transform 1 0 15202 0 1 -16552
box 70 126 186 240
use ptap  ptap_68
timestamp 1624298412
transform 1 0 17238 0 1 -16552
box 70 126 186 240
use ptap  ptap_67
timestamp 1624298412
transform 1 0 16220 0 1 -16552
box 70 126 186 240
use ptap  ptap_69
timestamp 1624298412
transform 1 0 18256 0 1 -16552
box 70 126 186 240
use ptap  ptap_70
timestamp 1624298412
transform 1 0 19274 0 1 -16552
box 70 126 186 240
use ptap  ptap_71
timestamp 1624298412
transform 1 0 20292 0 1 -16552
box 70 126 186 240
use ptap  ptap_72
timestamp 1624298412
transform 1 0 21310 0 1 -16552
box 70 126 186 240
use ptap  ptap_73
timestamp 1624298412
transform 1 0 22328 0 1 -16552
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_8
timestamp 1624298412
transform 1 0 12779 0 1 -15764
box -10209 -388 10209 388
use ptap  ptap_346
timestamp 1624298412
transform 1 0 -9296 0 1 -15858
box 70 126 186 240
use ptap  ptap_347
timestamp 1624298412
transform 1 0 -8278 0 1 -15858
box 70 126 186 240
use ptap  ptap_348
timestamp 1624298412
transform 1 0 -7260 0 1 -15858
box 70 126 186 240
use ptap  ptap_349
timestamp 1624298412
transform 1 0 -6242 0 1 -15858
box 70 126 186 240
use ptap  ptap_350
timestamp 1624298412
transform 1 0 -5224 0 1 -15858
box 70 126 186 240
use ptap  ptap_351
timestamp 1624298412
transform 1 0 -4206 0 1 -15858
box 70 126 186 240
use ptap  ptap_352
timestamp 1624298412
transform 1 0 -3188 0 1 -15858
box 70 126 186 240
use ptap  ptap_353
timestamp 1624298412
transform 1 0 -2170 0 1 -15858
box 70 126 186 240
use ptap  ptap_354
timestamp 1624298412
transform 1 0 -1152 0 1 -15858
box 70 126 186 240
use ptap  ptap_355
timestamp 1624298412
transform 1 0 -124 0 1 -15858
box 70 126 186 240
use ptap  ptap_54
timestamp 1624298412
transform 1 0 2998 0 1 -15316
box 70 126 186 240
use ptap  ptap_56
timestamp 1624298412
transform 1 0 5034 0 1 -15316
box 70 126 186 240
use ptap  ptap_55
timestamp 1624298412
transform 1 0 4016 0 1 -15316
box 70 126 186 240
use ptap  ptap_57
timestamp 1624298412
transform 1 0 6052 0 1 -15316
box 70 126 186 240
use ptap  ptap_58
timestamp 1624298412
transform 1 0 7070 0 1 -15316
box 70 126 186 240
use ptap  ptap_59
timestamp 1624298412
transform 1 0 8088 0 1 -15316
box 70 126 186 240
use ptap  ptap_40
timestamp 1624298412
transform 1 0 9106 0 1 -15316
box 70 126 186 240
use ptap  ptap_41
timestamp 1624298412
transform 1 0 10124 0 1 -15316
box 70 126 186 240
use ptap  ptap_42
timestamp 1624298412
transform 1 0 11142 0 1 -15316
box 70 126 186 240
use ptap  ptap_43
timestamp 1624298412
transform 1 0 12160 0 1 -15316
box 70 126 186 240
use ptap  ptap_44
timestamp 1624298412
transform 1 0 13178 0 1 -15316
box 70 126 186 240
use ptap  ptap_45
timestamp 1624298412
transform 1 0 14196 0 1 -15316
box 70 126 186 240
use ptap  ptap_46
timestamp 1624298412
transform 1 0 15214 0 1 -15316
box 70 126 186 240
use ptap  ptap_48
timestamp 1624298412
transform 1 0 17250 0 1 -15316
box 70 126 186 240
use ptap  ptap_47
timestamp 1624298412
transform 1 0 16232 0 1 -15316
box 70 126 186 240
use ptap  ptap_49
timestamp 1624298412
transform 1 0 18268 0 1 -15316
box 70 126 186 240
use ptap  ptap_50
timestamp 1624298412
transform 1 0 19286 0 1 -15316
box 70 126 186 240
use ptap  ptap_51
timestamp 1624298412
transform 1 0 20304 0 1 -15316
box 70 126 186 240
use ptap  ptap_52
timestamp 1624298412
transform 1 0 21322 0 1 -15316
box 70 126 186 240
use ptap  ptap_53
timestamp 1624298412
transform 1 0 22340 0 1 -15316
box 70 126 186 240
use ptap  ptap_356
timestamp 1624298412
transform 1 0 -9296 0 1 -15040
box 70 126 186 240
use ptap  ptap_357
timestamp 1624298412
transform 1 0 -8278 0 1 -15040
box 70 126 186 240
use ptap  ptap_358
timestamp 1624298412
transform 1 0 -7260 0 1 -15040
box 70 126 186 240
use ptap  ptap_360
timestamp 1624298412
transform 1 0 -5224 0 1 -15040
box 70 126 186 240
use ptap  ptap_359
timestamp 1624298412
transform 1 0 -6242 0 1 -15040
box 70 126 186 240
use ptap  ptap_361
timestamp 1624298412
transform 1 0 -4206 0 1 -15040
box 70 126 186 240
use ptap  ptap_363
timestamp 1624298412
transform 1 0 -2170 0 1 -15040
box 70 126 186 240
use ptap  ptap_362
timestamp 1624298412
transform 1 0 -3188 0 1 -15040
box 70 126 186 240
use ptap  ptap_364
timestamp 1624298412
transform 1 0 -1152 0 1 -15040
box 70 126 186 240
use ptap  ptap_365
timestamp 1624298412
transform 1 0 -124 0 1 -15040
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_MCKC3T  sky130_fd_pr__nfet_01v8_MCKC3T_7
timestamp 1624298412
transform 1 0 12779 0 1 -14532
box -10209 -388 10209 388
use ptap  ptap_366
timestamp 1624298412
transform 1 0 -9296 0 1 -14222
box 70 126 186 240
use ptap  ptap_368
timestamp 1624298412
transform 1 0 -7260 0 1 -14222
box 70 126 186 240
use ptap  ptap_367
timestamp 1624298412
transform 1 0 -8278 0 1 -14222
box 70 126 186 240
use ptap  ptap_369
timestamp 1624298412
transform 1 0 -6242 0 1 -14222
box 70 126 186 240
use ptap  ptap_370
timestamp 1624298412
transform 1 0 -5224 0 1 -14222
box 70 126 186 240
use ptap  ptap_371
timestamp 1624298412
transform 1 0 -4206 0 1 -14222
box 70 126 186 240
use ptap  ptap_372
timestamp 1624298412
transform 1 0 -3188 0 1 -14222
box 70 126 186 240
use ptap  ptap_373
timestamp 1624298412
transform 1 0 -2170 0 1 -14222
box 70 126 186 240
use ptap  ptap_374
timestamp 1624298412
transform 1 0 -1152 0 1 -14222
box 70 126 186 240
use ptap  ptap_375
timestamp 1624298412
transform 1 0 -124 0 1 -14222
box 70 126 186 240
use ptap  ptap_34
timestamp 1624298412
transform 1 0 3010 0 1 -14010
box 70 126 186 240
use ptap  ptap_36
timestamp 1624298412
transform 1 0 5046 0 1 -14010
box 70 126 186 240
use ptap  ptap_35
timestamp 1624298412
transform 1 0 4028 0 1 -14010
box 70 126 186 240
use ptap  ptap_37
timestamp 1624298412
transform 1 0 6064 0 1 -14010
box 70 126 186 240
use ptap  ptap_38
timestamp 1624298412
transform 1 0 7082 0 1 -14010
box 70 126 186 240
use ptap  ptap_39
timestamp 1624298412
transform 1 0 8100 0 1 -14010
box 70 126 186 240
use ptap  ptap_20
timestamp 1624298412
transform 1 0 9118 0 1 -14010
box 70 126 186 240
use ptap  ptap_21
timestamp 1624298412
transform 1 0 10136 0 1 -14010
box 70 126 186 240
use ptap  ptap_22
timestamp 1624298412
transform 1 0 11154 0 1 -14010
box 70 126 186 240
use ptap  ptap_23
timestamp 1624298412
transform 1 0 12172 0 1 -14010
box 70 126 186 240
use ptap  ptap_24
timestamp 1624298412
transform 1 0 13190 0 1 -14010
box 70 126 186 240
use ptap  ptap_25
timestamp 1624298412
transform 1 0 14208 0 1 -14010
box 70 126 186 240
use ptap  ptap_26
timestamp 1624298412
transform 1 0 15226 0 1 -14010
box 70 126 186 240
use ptap  ptap_28
timestamp 1624298412
transform 1 0 17262 0 1 -14010
box 70 126 186 240
use ptap  ptap_27
timestamp 1624298412
transform 1 0 16244 0 1 -14010
box 70 126 186 240
use ptap  ptap_29
timestamp 1624298412
transform 1 0 18280 0 1 -14010
box 70 126 186 240
use ptap  ptap_30
timestamp 1624298412
transform 1 0 19298 0 1 -14010
box 70 126 186 240
use ptap  ptap_31
timestamp 1624298412
transform 1 0 20316 0 1 -14010
box 70 126 186 240
use ptap  ptap_32
timestamp 1624298412
transform 1 0 21334 0 1 -14010
box 70 126 186 240
use ptap  ptap_33
timestamp 1624298412
transform 1 0 22352 0 1 -14010
box 70 126 186 240
use sky130_fd_pr__nfet_01v8_J5YDRX  sky130_fd_pr__nfet_01v8_J5YDRX_0
timestamp 1624298412
transform -1 0 12779 0 -1 -12745
box -10209 -797 10209 797
use sky130_fd_pr__nfet_01v8_lvt_XH9Q8F  sky130_fd_pr__nfet_01v8_lvt_XH9Q8F_0
timestamp 1624298412
transform 1 0 -4586 0 1 -14039
box -4610 -1615 4610 1615
use ptap  ptap_376
timestamp 1624298412
transform 1 0 -9296 0 1 -13404
box 70 126 186 240
use ptap  ptap_386
timestamp 1624298412
transform 1 0 -9296 0 1 -12586
box 70 126 186 240
use ptap  ptap_387
timestamp 1624298412
transform 1 0 -8278 0 1 -12586
box 70 126 186 240
use ptap  ptap_377
timestamp 1624298412
transform 1 0 -8278 0 1 -13404
box 70 126 186 240
use ptap  ptap_388
timestamp 1624298412
transform 1 0 -7260 0 1 -12586
box 70 126 186 240
use ptap  ptap_378
timestamp 1624298412
transform 1 0 -7260 0 1 -13404
box 70 126 186 240
use ptap  ptap_389
timestamp 1624298412
transform 1 0 -6242 0 1 -12586
box 70 126 186 240
use ptap  ptap_379
timestamp 1624298412
transform 1 0 -6242 0 1 -13404
box 70 126 186 240
use ptap  ptap_390
timestamp 1624298412
transform 1 0 -5224 0 1 -12586
box 70 126 186 240
use ptap  ptap_380
timestamp 1624298412
transform 1 0 -5224 0 1 -13404
box 70 126 186 240
use ptap  ptap_391
timestamp 1624298412
transform 1 0 -4206 0 1 -12586
box 70 126 186 240
use ptap  ptap_381
timestamp 1624298412
transform 1 0 -4206 0 1 -13404
box 70 126 186 240
use ptap  ptap_392
timestamp 1624298412
transform 1 0 -3188 0 1 -12586
box 70 126 186 240
use ptap  ptap_382
timestamp 1624298412
transform 1 0 -3188 0 1 -13404
box 70 126 186 240
use ptap  ptap_393
timestamp 1624298412
transform 1 0 -2170 0 1 -12586
box 70 126 186 240
use ptap  ptap_383
timestamp 1624298412
transform 1 0 -2170 0 1 -13404
box 70 126 186 240
use ptap  ptap_394
timestamp 1624298412
transform 1 0 -1152 0 1 -12586
box 70 126 186 240
use ptap  ptap_384
timestamp 1624298412
transform 1 0 -1152 0 1 -13404
box 70 126 186 240
use ptap  ptap_395
timestamp 1624298412
transform 1 0 -124 0 1 -12586
box 70 126 186 240
use ptap  ptap_385
timestamp 1624298412
transform 1 0 -124 0 1 -13404
box 70 126 186 240
use ptap  ptap_0
timestamp 1624298412
transform 1 0 2998 0 1 -11984
box 70 126 186 240
use ptap  ptap_1
timestamp 1624298412
transform 1 0 4016 0 1 -11984
box 70 126 186 240
use ptap  ptap_2
timestamp 1624298412
transform 1 0 5034 0 1 -11984
box 70 126 186 240
use ptap  ptap_3
timestamp 1624298412
transform 1 0 6052 0 1 -11984
box 70 126 186 240
use ptap  ptap_4
timestamp 1624298412
transform 1 0 7070 0 1 -11984
box 70 126 186 240
use ptap  ptap_5
timestamp 1624298412
transform 1 0 8088 0 1 -11984
box 70 126 186 240
use ptap  ptap_6
timestamp 1624298412
transform 1 0 9106 0 1 -11984
box 70 126 186 240
use ptap  ptap_7
timestamp 1624298412
transform 1 0 10124 0 1 -11984
box 70 126 186 240
use ptap  ptap_8
timestamp 1624298412
transform 1 0 11142 0 1 -11984
box 70 126 186 240
use ptap  ptap_9
timestamp 1624298412
transform 1 0 12160 0 1 -11984
box 70 126 186 240
use ptap  ptap_10
timestamp 1624298412
transform 1 0 13178 0 1 -11984
box 70 126 186 240
use ptap  ptap_11
timestamp 1624298412
transform 1 0 14196 0 1 -11984
box 70 126 186 240
use ptap  ptap_12
timestamp 1624298412
transform 1 0 15214 0 1 -11984
box 70 126 186 240
use ptap  ptap_13
timestamp 1624298412
transform 1 0 16232 0 1 -11984
box 70 126 186 240
use ptap  ptap_14
timestamp 1624298412
transform 1 0 17250 0 1 -11984
box 70 126 186 240
use ptap  ptap_15
timestamp 1624298412
transform 1 0 18268 0 1 -11984
box 70 126 186 240
use ptap  ptap_16
timestamp 1624298412
transform 1 0 19286 0 1 -11984
box 70 126 186 240
use ptap  ptap_17
timestamp 1624298412
transform 1 0 20304 0 1 -11984
box 70 126 186 240
use ptap  ptap_18
timestamp 1624298412
transform 1 0 21322 0 1 -11984
box 70 126 186 240
use ptap  ptap_19
timestamp 1624298412
transform 1 0 22340 0 1 -11984
box 70 126 186 240
use ntap  ntap_162 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/ntap
timestamp 1624298412
transform 1 0 2348 0 1 -9532
box 250 218 480 436
use ntap  ntap_161
timestamp 1624298412
transform 1 0 3366 0 1 -9532
box 250 218 480 436
use ntap  ntap_160
timestamp 1624298412
transform 1 0 4384 0 1 -9532
box 250 218 480 436
use ntap  ntap_159
timestamp 1624298412
transform 1 0 5402 0 1 -9532
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_3
timestamp 1624298412
transform 1 0 15126 0 1 -9140
box -7700 -400 7700 400
use sky130_fd_pr__pfet_01v8_lvt_DHLX6D  sky130_fd_pr__pfet_01v8_lvt_DHLX6D_3
timestamp 1624298412
transform 1 0 4223 0 1 -8572
box -2101 -400 2101 400
use ntap  ntap_122
timestamp 1624298412
transform 1 0 6924 0 1 -8820
box 250 218 480 436
use ntap  ntap_123
timestamp 1624298412
transform 1 0 7942 0 1 -8820
box 250 218 480 436
use ntap  ntap_124
timestamp 1624298412
transform 1 0 8960 0 1 -8820
box 250 218 480 436
use ntap  ntap_125
timestamp 1624298412
transform 1 0 9978 0 1 -8820
box 250 218 480 436
use ntap  ntap_126
timestamp 1624298412
transform 1 0 10996 0 1 -8820
box 250 218 480 436
use ntap  ntap_127
timestamp 1624298412
transform 1 0 12014 0 1 -8820
box 250 218 480 436
use ntap  ntap_113
timestamp 1624298412
transform 1 0 14050 0 1 -8820
box 250 218 480 436
use ntap  ntap_112
timestamp 1624298412
transform 1 0 13032 0 1 -8820
box 250 218 480 436
use ntap  ntap_114
timestamp 1624298412
transform 1 0 15068 0 1 -8820
box 250 218 480 436
use ntap  ntap_115
timestamp 1624298412
transform 1 0 16086 0 1 -8820
box 250 218 480 436
use ntap  ntap_116
timestamp 1624298412
transform 1 0 17104 0 1 -8820
box 250 218 480 436
use ntap  ntap_117
timestamp 1624298412
transform 1 0 18122 0 1 -8820
box 250 218 480 436
use ntap  ntap_118
timestamp 1624298412
transform 1 0 19140 0 1 -8820
box 250 218 480 436
use ntap  ntap_119
timestamp 1624298412
transform 1 0 20158 0 1 -8820
box 250 218 480 436
use ntap  ntap_120
timestamp 1624298412
transform 1 0 21176 0 1 -8820
box 250 218 480 436
use ntap  ntap_121
timestamp 1624298412
transform 1 0 22194 0 1 -8820
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_DHLX6D  sky130_fd_pr__pfet_01v8_lvt_DHLX6D_2
timestamp 1624298412
transform 1 0 4223 0 1 -7540
box -2101 -400 2101 400
use ntap  ntap_156
timestamp 1624298412
transform 1 0 3860 0 1 -8380
box 250 218 480 436
use ntap  ntap_157
timestamp 1624298412
transform 1 0 2842 0 1 -8380
box 250 218 480 436
use ntap  ntap_158
timestamp 1624298412
transform 1 0 1824 0 1 -8380
box 250 218 480 436
use ntap  ntap_155
timestamp 1624298412
transform 1 0 4878 0 1 -8380
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_2
timestamp 1624298412
transform 1 0 15126 0 1 -7884
box -7700 -400 7700 400
use sky130_fd_pr__pfet_01v8_lvt_DHLX6D  sky130_fd_pr__pfet_01v8_lvt_DHLX6D_1
timestamp 1624298412
transform 1 0 4223 0 1 -6508
box -2101 -400 2101 400
use ntap  ntap_154
timestamp 1624298412
transform 1 0 1834 0 1 -7352
box 250 218 480 436
use ntap  ntap_153
timestamp 1624298412
transform 1 0 2852 0 1 -7352
box 250 218 480 436
use ntap  ntap_152
timestamp 1624298412
transform 1 0 3870 0 1 -7352
box 250 218 480 436
use ntap  ntap_106
timestamp 1624298412
transform 1 0 7060 0 1 -7576
box 250 218 480 436
use ntap  ntap_107
timestamp 1624298412
transform 1 0 8078 0 1 -7576
box 250 218 480 436
use ntap  ntap_108
timestamp 1624298412
transform 1 0 9096 0 1 -7576
box 250 218 480 436
use ntap  ntap_109
timestamp 1624298412
transform 1 0 10114 0 1 -7576
box 250 218 480 436
use ntap  ntap_110
timestamp 1624298412
transform 1 0 11132 0 1 -7576
box 250 218 480 436
use ntap  ntap_111
timestamp 1624298412
transform 1 0 12150 0 1 -7576
box 250 218 480 436
use ntap  ntap_96
timestamp 1624298412
transform 1 0 13168 0 1 -7576
box 250 218 480 436
use ntap  ntap_97
timestamp 1624298412
transform 1 0 14186 0 1 -7576
box 250 218 480 436
use ntap  ntap_98
timestamp 1624298412
transform 1 0 15204 0 1 -7576
box 250 218 480 436
use ntap  ntap_99
timestamp 1624298412
transform 1 0 16222 0 1 -7576
box 250 218 480 436
use ntap  ntap_100
timestamp 1624298412
transform 1 0 17240 0 1 -7576
box 250 218 480 436
use ntap  ntap_101
timestamp 1624298412
transform 1 0 18258 0 1 -7576
box 250 218 480 436
use ntap  ntap_102
timestamp 1624298412
transform 1 0 19276 0 1 -7576
box 250 218 480 436
use ntap  ntap_151
timestamp 1624298412
transform 1 0 4888 0 1 -7352
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_0
timestamp 1624298412
transform 1 0 15126 0 1 -6628
box -7700 -400 7700 400
use ntap  ntap_103
timestamp 1624298412
transform 1 0 20294 0 1 -7576
box 250 218 480 436
use ntap  ntap_104
timestamp 1624298412
transform 1 0 21312 0 1 -7576
box 250 218 480 436
use ntap  ntap_105
timestamp 1624298412
transform 1 0 22330 0 1 -7576
box 250 218 480 436
use ntap  ntap_149
timestamp 1624298412
transform 1 0 2842 0 1 -6324
box 250 218 480 436
use ntap  ntap_150
timestamp 1624298412
transform 1 0 1824 0 1 -6324
box 250 218 480 436
use ntap  ntap_148
timestamp 1624298412
transform 1 0 3860 0 1 -6324
box 250 218 480 436
use ntap  ntap_147
timestamp 1624298412
transform 1 0 4878 0 1 -6324
box 250 218 480 436
use ntap  ntap_90
timestamp 1624298412
transform 1 0 7036 0 1 -6308
box 250 218 480 436
use ntap  ntap_91
timestamp 1624298412
transform 1 0 8054 0 1 -6308
box 250 218 480 436
use ntap  ntap_93
timestamp 1624298412
transform 1 0 10090 0 1 -6308
box 250 218 480 436
use ntap  ntap_92
timestamp 1624298412
transform 1 0 9072 0 1 -6308
box 250 218 480 436
use ntap  ntap_94
timestamp 1624298412
transform 1 0 11108 0 1 -6308
box 250 218 480 436
use ntap  ntap_95
timestamp 1624298412
transform 1 0 12126 0 1 -6308
box 250 218 480 436
use ntap  ntap_80
timestamp 1624298412
transform 1 0 13144 0 1 -6308
box 250 218 480 436
use ntap  ntap_81
timestamp 1624298412
transform 1 0 14162 0 1 -6308
box 250 218 480 436
use ntap  ntap_82
timestamp 1624298412
transform 1 0 15180 0 1 -6308
box 250 218 480 436
use ntap  ntap_83
timestamp 1624298412
transform 1 0 16198 0 1 -6308
box 250 218 480 436
use ntap  ntap_84
timestamp 1624298412
transform 1 0 17216 0 1 -6308
box 250 218 480 436
use ntap  ntap_85
timestamp 1624298412
transform 1 0 18234 0 1 -6308
box 250 218 480 436
use ntap  ntap_86
timestamp 1624298412
transform 1 0 19252 0 1 -6308
box 250 218 480 436
use ntap  ntap_87
timestamp 1624298412
transform 1 0 20270 0 1 -6308
box 250 218 480 436
use ntap  ntap_89
timestamp 1624298412
transform 1 0 22306 0 1 -6308
box 250 218 480 436
use ntap  ntap_88
timestamp 1624298412
transform 1 0 21288 0 1 -6308
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_DHLX6D  sky130_fd_pr__pfet_01v8_lvt_DHLX6D_0
timestamp 1624298412
transform 1 0 4223 0 1 -5476
box -2101 -400 2101 400
use sky130_fd_pr__pfet_01v8_MSJKJ2  sky130_fd_pr__pfet_01v8_MSJKJ2_1
timestamp 1624298412
transform 1 0 15126 0 1 -5372
box -7700 -400 7700 400
use ntap  ntap_146
timestamp 1624298412
transform 1 0 2348 0 1 -5170
box 250 218 480 436
use ntap  ntap_145
timestamp 1624298412
transform 1 0 3366 0 1 -5170
box 250 218 480 436
use ntap  ntap_144
timestamp 1624298412
transform 1 0 4384 0 1 -5170
box 250 218 480 436
use ntap  ntap_143
timestamp 1624298412
transform 1 0 5402 0 1 -5170
box 250 218 480 436
use ntap  ntap_74
timestamp 1624298412
transform 1 0 6946 0 1 -4860
box 250 218 480 436
use ntap  ntap_75
timestamp 1624298412
transform 1 0 7964 0 1 -4860
box 250 218 480 436
use ntap  ntap_76
timestamp 1624298412
transform 1 0 8982 0 1 -4860
box 250 218 480 436
use ntap  ntap_77
timestamp 1624298412
transform 1 0 10000 0 1 -4860
box 250 218 480 436
use ntap  ntap_78
timestamp 1624298412
transform 1 0 11018 0 1 -4860
box 250 218 480 436
use ntap  ntap_79
timestamp 1624298412
transform 1 0 12036 0 1 -4860
box 250 218 480 436
use ntap  ntap_64
timestamp 1624298412
transform 1 0 13054 0 1 -4860
box 250 218 480 436
use ntap  ntap_65
timestamp 1624298412
transform 1 0 14072 0 1 -4860
box 250 218 480 436
use ntap  ntap_66
timestamp 1624298412
transform 1 0 15090 0 1 -4860
box 250 218 480 436
use ntap  ntap_67
timestamp 1624298412
transform 1 0 16108 0 1 -4860
box 250 218 480 436
use ntap  ntap_68
timestamp 1624298412
transform 1 0 17126 0 1 -4860
box 250 218 480 436
use ntap  ntap_69
timestamp 1624298412
transform 1 0 18144 0 1 -4860
box 250 218 480 436
use ntap  ntap_70
timestamp 1624298412
transform 1 0 19162 0 1 -4860
box 250 218 480 436
use ntap  ntap_71
timestamp 1624298412
transform 1 0 20180 0 1 -4860
box 250 218 480 436
use ntap  ntap_72
timestamp 1624298412
transform 1 0 21198 0 1 -4860
box 250 218 480 436
use ntap  ntap_73
timestamp 1624298412
transform 1 0 22216 0 1 -4860
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_SH2KEA  sky130_fd_pr__pfet_01v8_lvt_SH2KEA_1
timestamp 1624298412
transform 1 0 14825 0 1 -3768
box -7191 -400 7191 400
use ntap  ntap_142
timestamp 1624298412
transform 1 0 7340 0 1 -3582
box 250 218 480 436
use ntap  ntap_141
timestamp 1624298412
transform 1 0 8358 0 1 -3582
box 250 218 480 436
use ntap  ntap_140
timestamp 1624298412
transform 1 0 9376 0 1 -3582
box 250 218 480 436
use ntap  ntap_139
timestamp 1624298412
transform 1 0 10394 0 1 -3582
box 250 218 480 436
use ntap  ntap_138
timestamp 1624298412
transform 1 0 11412 0 1 -3582
box 250 218 480 436
use ntap  ntap_137
timestamp 1624298412
transform 1 0 12430 0 1 -3582
box 250 218 480 436
use ntap  ntap_136
timestamp 1624298412
transform 1 0 13448 0 1 -3582
box 250 218 480 436
use ntap  ntap_135
timestamp 1624298412
transform 1 0 14466 0 1 -3582
box 250 218 480 436
use ntap  ntap_134
timestamp 1624298412
transform 1 0 15484 0 1 -3582
box 250 218 480 436
use ntap  ntap_133
timestamp 1624298412
transform 1 0 16502 0 1 -3582
box 250 218 480 436
use ntap  ntap_132
timestamp 1624298412
transform 1 0 17520 0 1 -3582
box 250 218 480 436
use ntap  ntap_131
timestamp 1624298412
transform 1 0 18538 0 1 -3582
box 250 218 480 436
use ntap  ntap_130
timestamp 1624298412
transform 1 0 19556 0 1 -3582
box 250 218 480 436
use ntap  ntap_128
timestamp 1624298412
transform 1 0 20574 0 1 -3582
box 250 218 480 436
use ntap  ntap_129
timestamp 1624298412
transform 1 0 21592 0 1 -3582
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_SH2KEA  sky130_fd_pr__pfet_01v8_lvt_SH2KEA_0
timestamp 1624298412
transform 1 0 14825 0 1 -2736
box -7191 -400 7191 400
use ntap  ntap_58
timestamp 1624298412
transform 1 0 6652 0 1 -2234
box 250 218 480 436
use ntap  ntap_59
timestamp 1624298412
transform 1 0 7670 0 1 -2234
box 250 218 480 436
use ntap  ntap_60
timestamp 1624298412
transform 1 0 8688 0 1 -2234
box 250 218 480 436
use ntap  ntap_61
timestamp 1624298412
transform 1 0 9706 0 1 -2234
box 250 218 480 436
use ntap  ntap_62
timestamp 1624298412
transform 1 0 10724 0 1 -2234
box 250 218 480 436
use ntap  ntap_63
timestamp 1624298412
transform 1 0 11742 0 1 -2234
box 250 218 480 436
use ntap  ntap_48
timestamp 1624298412
transform 1 0 12760 0 1 -2234
box 250 218 480 436
use ntap  ntap_49
timestamp 1624298412
transform 1 0 13778 0 1 -2234
box 250 218 480 436
use ntap  ntap_50
timestamp 1624298412
transform 1 0 14796 0 1 -2234
box 250 218 480 436
use ntap  ntap_51
timestamp 1624298412
transform 1 0 15814 0 1 -2234
box 250 218 480 436
use ntap  ntap_52
timestamp 1624298412
transform 1 0 16832 0 1 -2234
box 250 218 480 436
use ntap  ntap_53
timestamp 1624298412
transform 1 0 17850 0 1 -2234
box 250 218 480 436
use ntap  ntap_54
timestamp 1624298412
transform 1 0 18868 0 1 -2234
box 250 218 480 436
use ntap  ntap_55
timestamp 1624298412
transform 1 0 19886 0 1 -2234
box 250 218 480 436
use ntap  ntap_56
timestamp 1624298412
transform 1 0 20904 0 1 -2234
box 250 218 480 436
use ntap  ntap_57
timestamp 1624298412
transform 1 0 21922 0 1 -2234
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_2
timestamp 1624298412
transform 1 0 14649 0 1 -1098
box -8209 -400 8209 400
use ntap  ntap_42
timestamp 1624298412
transform 1 0 6652 0 1 -852
box 250 218 480 436
use ntap  ntap_43
timestamp 1624298412
transform 1 0 7670 0 1 -852
box 250 218 480 436
use ntap  ntap_44
timestamp 1624298412
transform 1 0 8688 0 1 -852
box 250 218 480 436
use ntap  ntap_45
timestamp 1624298412
transform 1 0 9706 0 1 -852
box 250 218 480 436
use ntap  ntap_46
timestamp 1624298412
transform 1 0 10724 0 1 -852
box 250 218 480 436
use ntap  ntap_47
timestamp 1624298412
transform 1 0 11742 0 1 -852
box 250 218 480 436
use ntap  ntap_32
timestamp 1624298412
transform 1 0 12760 0 1 -852
box 250 218 480 436
use ntap  ntap_33
timestamp 1624298412
transform 1 0 13778 0 1 -852
box 250 218 480 436
use ntap  ntap_34
timestamp 1624298412
transform 1 0 14796 0 1 -852
box 250 218 480 436
use ntap  ntap_35
timestamp 1624298412
transform 1 0 15814 0 1 -852
box 250 218 480 436
use ntap  ntap_36
timestamp 1624298412
transform 1 0 16832 0 1 -852
box 250 218 480 436
use ntap  ntap_37
timestamp 1624298412
transform 1 0 17850 0 1 -852
box 250 218 480 436
use ntap  ntap_38
timestamp 1624298412
transform 1 0 18868 0 1 -852
box 250 218 480 436
use ntap  ntap_39
timestamp 1624298412
transform 1 0 19886 0 1 -852
box 250 218 480 436
use ntap  ntap_40
timestamp 1624298412
transform 1 0 20904 0 1 -852
box 250 218 480 436
use ntap  ntap_41
timestamp 1624298412
transform 1 0 21922 0 1 -852
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_1
timestamp 1624298412
transform 1 0 14649 0 1 38
box -8209 -400 8209 400
use ntap  ntap_26
timestamp 1624298412
transform 1 0 6674 0 1 280
box 250 218 480 436
use ntap  ntap_27
timestamp 1624298412
transform 1 0 7692 0 1 280
box 250 218 480 436
use ntap  ntap_28
timestamp 1624298412
transform 1 0 8710 0 1 280
box 250 218 480 436
use ntap  ntap_29
timestamp 1624298412
transform 1 0 9728 0 1 280
box 250 218 480 436
use ntap  ntap_30
timestamp 1624298412
transform 1 0 10746 0 1 280
box 250 218 480 436
use ntap  ntap_31
timestamp 1624298412
transform 1 0 11764 0 1 280
box 250 218 480 436
use ntap  ntap_16
timestamp 1624298412
transform 1 0 12782 0 1 280
box 250 218 480 436
use ntap  ntap_17
timestamp 1624298412
transform 1 0 13800 0 1 280
box 250 218 480 436
use ntap  ntap_18
timestamp 1624298412
transform 1 0 14818 0 1 280
box 250 218 480 436
use ntap  ntap_19
timestamp 1624298412
transform 1 0 15836 0 1 280
box 250 218 480 436
use ntap  ntap_20
timestamp 1624298412
transform 1 0 16854 0 1 280
box 250 218 480 436
use ntap  ntap_21
timestamp 1624298412
transform 1 0 17872 0 1 280
box 250 218 480 436
use ntap  ntap_22
timestamp 1624298412
transform 1 0 18890 0 1 280
box 250 218 480 436
use ntap  ntap_23
timestamp 1624298412
transform 1 0 19908 0 1 280
box 250 218 480 436
use ntap  ntap_24
timestamp 1624298412
transform 1 0 20926 0 1 280
box 250 218 480 436
use ntap  ntap_25
timestamp 1624298412
transform 1 0 21944 0 1 280
box 250 218 480 436
use sky130_fd_pr__pfet_01v8_lvt_V2JKJ2  sky130_fd_pr__pfet_01v8_lvt_V2JKJ2_0
timestamp 1624298412
transform 1 0 14649 0 1 1174
box -8209 -400 8209 400
use ntap  ntap_0
timestamp 1624298412
transform 1 0 6652 0 1 1434
box 250 218 480 436
use ntap  ntap_1
timestamp 1624298412
transform 1 0 7670 0 1 1434
box 250 218 480 436
use ntap  ntap_2
timestamp 1624298412
transform 1 0 8688 0 1 1434
box 250 218 480 436
use ntap  ntap_3
timestamp 1624298412
transform 1 0 9706 0 1 1434
box 250 218 480 436
use ntap  ntap_4
timestamp 1624298412
transform 1 0 10724 0 1 1434
box 250 218 480 436
use ntap  ntap_5
timestamp 1624298412
transform 1 0 11742 0 1 1434
box 250 218 480 436
use ntap  ntap_6
timestamp 1624298412
transform 1 0 12760 0 1 1434
box 250 218 480 436
use ntap  ntap_7
timestamp 1624298412
transform 1 0 13778 0 1 1434
box 250 218 480 436
use ntap  ntap_8
timestamp 1624298412
transform 1 0 14796 0 1 1434
box 250 218 480 436
use ntap  ntap_9
timestamp 1624298412
transform 1 0 15814 0 1 1434
box 250 218 480 436
use ntap  ntap_10
timestamp 1624298412
transform 1 0 16832 0 1 1434
box 250 218 480 436
use ntap  ntap_11
timestamp 1624298412
transform 1 0 17850 0 1 1434
box 250 218 480 436
use ntap  ntap_12
timestamp 1624298412
transform 1 0 18868 0 1 1434
box 250 218 480 436
use ntap  ntap_13
timestamp 1624298412
transform 1 0 19886 0 1 1434
box 250 218 480 436
use ntap  ntap_14
timestamp 1624298412
transform 1 0 20904 0 1 1434
box 250 218 480 436
use ntap  ntap_15
timestamp 1624298412
transform 1 0 21922 0 1 1434
box 250 218 480 436
<< labels >>
flabel metal1 -8078 -12352 -8078 -12352 1 FreeSans 480 0 0 0 vbias1
flabel metal1 -6206 -19026 -6206 -19026 1 FreeSans 480 0 0 0 vbias2
flabel metal1 23180 -19318 23204 -19288 1 FreeSans 480 0 0 0 VSS
flabel metal1 23556 -18470 23556 -18470 1 FreeSans 480 0 0 0 vbias3
flabel metal1 23300 -18264 23300 -18264 1 FreeSans 480 0 0 0 vcascnm
flabel metal1 23436 -22496 23436 -22496 1 FreeSans 480 0 0 0 vbias4
flabel metal1 2138 -18102 2166 -18072 1 FreeSans 480 0 0 0 vtail_cascn
flabel metal1 2456 -14760 2488 -14720 1 FreeSans 480 0 0 0 vcascnp
flabel metal1 3322 -11898 3412 -11868 1 FreeSans 480 0 0 0 M8d
flabel metal1 2244 -18362 2282 -18326 1 FreeSans 480 0 0 0 vmirror
flabel metal1 22938 -16630 22974 -16600 1 FreeSans 480 0 0 0 M16d
flabel metal1 -10646 -21540 -10618 -21496 1 FreeSans 480 0 0 0 vip
flabel metal1 954 -21536 986 -21498 1 FreeSans 480 0 0 0 vim
flabel metal1 -5202 -24966 -5106 -24930 1 FreeSans 480 0 0 0 ibiasn
flabel metal1 -52 -22240 -4 -22216 1 FreeSans 480 0 0 0 vtail_cascn
flabel metal4 -10920 -26744 -10894 -26722 1 FreeSans 3200 0 0 0 VSS
flabel metal2 -6564 -19934 -6516 -19918 1 FreeSans 480 0 0 0 vcascpp
flabel metal1 -9488 -22168 -9456 -22140 1 FreeSans 480 0 0 0 vcascpm
flabel metal4 -11704 3910 -11678 4004 1 FreeSans 3200 0 0 0 VDD
flabel metal4 594 -11002 614 -10982 1 FreeSans 480 0 0 0 vo
flabel metal1 22608 -8372 22614 -8354 1 FreeSans 480 0 0 0 vo
flabel metal1 7498 -1550 7530 -1518 1 FreeSans 480 0 0 0 M9d
flabel metal1 2932 -5008 3004 -4978 1 FreeSans 480 0 0 0 vcascnm
flabel metal1 5656 -5000 5698 -4978 1 FreeSans 480 0 0 0 vcascnp
flabel metal1 4210 -5038 4236 -5000 1 FreeSans 480 0 0 0 vtail_cascp
flabel metal1 3698 -9046 3728 -9020 1 FreeSans 480 0 0 0 vip
flabel metal1 4706 -9050 4736 -9016 1 FreeSans 480 0 0 0 vim
flabel metal2 20172 -4390 20234 -4362 1 FreeSans 480 0 0 0 vmirror
flabel metal1 16210 -2186 16262 -2160 1 FreeSans 480 0 0 0 VDD
flabel metal2 10446 -3228 10514 -3198 1 FreeSans 480 0 0 0 vcascpp
flabel metal2 10670 -4260 10722 -4226 1 FreeSans 480 0 0 0 vcascpm
flabel metal2 8324 1884 8324 1884 1 FreeSans 480 0 0 0 vbias1
flabel metal2 9302 1622 9332 1650 1 FreeSans 480 0 0 0 VDD
flabel metal1 6346 610 6380 632 1 FreeSans 480 0 0 0 M7d
flabel metal2 7734 486 7792 522 1 FreeSans 480 0 0 0 M13d
flabel metal2 9760 -1694 9838 -1660 1 FreeSans 480 0 0 0 vtail_cascp
flabel metal1 17510 -5860 17546 -5832 1 FreeSans 480 0 0 0 VDD
flabel metal2 11866 -9908 11920 -9874 1 FreeSans 480 0 0 0 M8d
flabel metal2 12290 -4920 12372 -4888 1 FreeSans 480 0 0 0 vbias2
flabel metal2 16840 -7430 16902 -7400 1 FreeSans 480 0 0 0 M16d
flabel metal2 16432 -7118 16496 -7086 1 FreeSans 480 0 0 0 M13d
flabel metal1 7324 -5080 7364 -5046 1 FreeSans 480 0 0 0 M7d
flabel metal2 22394 -7218 22456 -7186 1 FreeSans 480 0 0 0 vmirror
flabel metal2 20508 -7328 20558 -7292 1 FreeSans 480 0 0 0 vcascpm
flabel metal2 20560 -8376 20652 -8344 1 FreeSans 480 0 0 0 vcascpp
flabel metal2 7618 -6048 7618 -6048 1 FreeSans 480 0 0 0 vbias1
flabel metal2 7488 -9634 7544 -9600 1 FreeSans 480 0 0 0 M9d
<< properties >>
string FIXED_BBOX -10872 -26372 24872 -10428
<< end >>

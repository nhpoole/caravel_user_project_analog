magic
tech sky130A
timestamp 1624300568
<< viali >>
rect 2052 206 2076 230
rect 144 144 168 168
rect 260 164 284 188
rect 1137 168 1161 192
rect 390 122 414 146
rect 2013 142 2037 166
rect 2099 142 2123 166
rect 2170 144 2194 168
rect 2221 142 2245 166
rect 192 97 216 121
rect 1263 116 1287 140
rect 943 91 967 115
rect 1817 91 1841 115
rect 1093 -39 1117 -15
rect 390 -63 414 -39
rect 1818 -41 1842 -17
rect 1263 -66 1287 -42
rect 260 -93 284 -69
rect 1140 -95 1164 -71
<< metal1 >>
rect -5 332 43 335
rect 43 284 66 332
rect -5 281 43 284
rect -36 203 257 233
rect 287 203 290 233
rect 2046 230 2197 233
rect 2046 206 2052 230
rect 2076 206 2197 230
rect 2046 203 2197 206
rect 257 188 287 203
rect 1134 195 1164 198
rect -36 168 174 171
rect -36 144 144 168
rect 168 144 174 168
rect 257 164 260 188
rect 284 164 287 188
rect 1131 165 1134 195
rect 1164 165 1167 195
rect 2096 169 2126 172
rect 1967 166 2043 169
rect 257 158 287 164
rect 1134 162 1164 165
rect -36 141 174 144
rect 387 146 417 152
rect 387 124 390 146
rect 186 122 390 124
rect 414 122 417 146
rect 186 121 417 122
rect 186 97 192 121
rect 216 97 417 121
rect 1260 140 1290 146
rect 1260 118 1263 140
rect 186 94 417 97
rect 937 116 1263 118
rect 1287 116 1290 140
rect 1967 142 2013 166
rect 2037 142 2043 166
rect 1967 139 2043 142
rect 2093 139 2096 169
rect 2126 139 2129 169
rect 2167 168 2197 203
rect 2167 144 2170 168
rect 2194 144 2197 168
rect 1812 118 1842 121
rect 1967 118 1997 139
rect 2096 136 2126 139
rect 2167 138 2197 144
rect 2215 166 2344 169
rect 2215 142 2221 166
rect 2245 142 2344 166
rect 2215 139 2344 142
rect 937 115 1290 116
rect 937 91 943 115
rect 967 91 1290 115
rect 937 88 1290 91
rect 1811 88 1812 118
rect 1842 88 1997 118
rect 1812 85 1842 88
rect -5 12 116 60
rect 1087 -15 1290 -12
rect 1967 -14 1997 -11
rect 387 -36 417 -33
rect 257 -66 287 -63
rect 384 -66 387 -36
rect 417 -66 420 -36
rect 1087 -39 1093 -15
rect 1117 -39 1290 -15
rect 1087 -42 1290 -39
rect 254 -96 257 -66
rect 287 -96 290 -66
rect 387 -69 417 -66
rect 1137 -68 1167 -65
rect 1260 -66 1263 -42
rect 1287 -66 1290 -42
rect 1812 -17 1967 -14
rect 1812 -41 1818 -17
rect 1842 -41 1967 -17
rect 1812 -44 1967 -41
rect 1967 -47 1997 -44
rect 257 -99 287 -96
rect 1134 -98 1137 -68
rect 1167 -98 1170 -68
rect 1260 -72 1290 -66
rect 1137 -101 1167 -98
rect -5 -212 43 -209
rect 43 -260 240 -212
rect -5 -263 43 -260
<< via1 >>
rect -5 284 43 332
rect 257 203 287 233
rect 1134 192 1164 195
rect 1134 168 1137 192
rect 1137 168 1161 192
rect 1161 168 1164 192
rect 1134 165 1164 168
rect 2096 166 2126 169
rect 2096 142 2099 166
rect 2099 142 2123 166
rect 2123 142 2126 166
rect 2096 139 2126 142
rect 1812 115 1842 118
rect 1812 91 1817 115
rect 1817 91 1841 115
rect 1841 91 1842 115
rect 1812 88 1842 91
rect 387 -39 417 -36
rect 387 -63 390 -39
rect 390 -63 414 -39
rect 414 -63 417 -39
rect 387 -66 417 -63
rect 257 -69 287 -66
rect 257 -93 260 -69
rect 260 -93 284 -69
rect 284 -93 287 -69
rect 257 -96 287 -93
rect 1967 -44 1997 -14
rect 1137 -71 1167 -68
rect 1137 -95 1140 -71
rect 1140 -95 1164 -71
rect 1164 -95 1167 -71
rect 1137 -98 1167 -95
rect -5 -260 43 -212
<< metal2 >>
rect -8 284 -5 332
rect 43 284 46 332
rect -5 -212 43 284
rect 257 233 287 236
rect 255 203 257 233
rect 287 203 1166 233
rect 257 -66 287 203
rect 1134 195 1164 203
rect 1134 162 1164 165
rect 1967 139 2096 169
rect 2126 139 2129 169
rect 1809 88 1812 118
rect 1842 88 1845 118
rect 1812 51 1842 88
rect 387 21 1842 51
rect 387 -36 417 21
rect 1967 -14 1997 139
rect 1964 -44 1967 -14
rect 1997 -44 2000 -14
rect 387 -69 417 -66
rect 1137 -68 1167 -65
rect 257 -107 287 -96
rect 1137 -107 1167 -98
rect 257 -137 1167 -107
rect -8 -260 -5 -212
rect 43 -260 46 -212
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624298412
transform 1 0 250 0 1 36
box -19 -24 893 296
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1624298412
transform 1 0 250 0 -1 36
box -19 -24 893 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624298412
transform 1 0 204 0 -1 36
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1624298412
transform 1 0 66 0 1 36
box -19 -24 65 296
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624299007
transform 1 0 112 0 1 36
box -19 -24 157 296
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1624298412
transform 1 0 1124 0 1 36
box -19 -24 893 296
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1624298412
transform 1 0 1124 0 -1 36
box -19 -24 893 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1624298412
transform 1 0 1998 0 -1 36
box -19 -24 65 296
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1624298412
transform 1 0 2274 0 1 36
box -19 -24 65 296
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1624299007
transform 1 0 2136 0 1 36
box -19 -24 157 296
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624299007
transform -1 0 2136 0 1 36
box -19 -24 157 296
<< labels >>
flabel metal2 10 251 13 253 1 FreeSans 240 0 0 0 VDD
flabel metal1 47 50 48 52 1 FreeSans 240 0 0 0 VSS
flabel metal1 -26 155 -22 159 1 FreeSans 240 0 0 0 trigb
flabel metal1 -26 217 -21 221 1 FreeSans 240 0 0 0 clk
flabel metal1 2322 152 2325 154 1 FreeSans 240 0 0 0 pulse
<< end >>

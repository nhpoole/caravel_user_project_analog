magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nwell >>
rect -1439 -200 1439 200
<< pmos >>
rect -1345 -100 -945 100
rect -887 -100 -487 100
rect -429 -100 -29 100
rect 29 -100 429 100
rect 487 -100 887 100
rect 945 -100 1345 100
<< pdiff >>
rect -1403 88 -1345 100
rect -1403 -88 -1391 88
rect -1357 -88 -1345 88
rect -1403 -100 -1345 -88
rect -945 88 -887 100
rect -945 -88 -933 88
rect -899 -88 -887 88
rect -945 -100 -887 -88
rect -487 88 -429 100
rect -487 -88 -475 88
rect -441 -88 -429 88
rect -487 -100 -429 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 429 88 487 100
rect 429 -88 441 88
rect 475 -88 487 88
rect 429 -100 487 -88
rect 887 88 945 100
rect 887 -88 899 88
rect 933 -88 945 88
rect 887 -100 945 -88
rect 1345 88 1403 100
rect 1345 -88 1357 88
rect 1391 -88 1403 88
rect 1345 -100 1403 -88
<< pdiffc >>
rect -1391 -88 -1357 88
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect 1357 -88 1391 88
<< poly >>
rect -1271 181 -1019 197
rect -1271 164 -1255 181
rect -1345 147 -1255 164
rect -1035 164 -1019 181
rect -813 181 -561 197
rect -813 164 -797 181
rect -1035 147 -945 164
rect -1345 100 -945 147
rect -887 147 -797 164
rect -577 164 -561 181
rect -355 181 -103 197
rect -355 164 -339 181
rect -577 147 -487 164
rect -887 100 -487 147
rect -429 147 -339 164
rect -119 164 -103 181
rect 103 181 355 197
rect 103 164 119 181
rect -119 147 -29 164
rect -429 100 -29 147
rect 29 147 119 164
rect 339 164 355 181
rect 561 181 813 197
rect 561 164 577 181
rect 339 147 429 164
rect 29 100 429 147
rect 487 147 577 164
rect 797 164 813 181
rect 1019 181 1271 197
rect 1019 164 1035 181
rect 797 147 887 164
rect 487 100 887 147
rect 945 147 1035 164
rect 1255 164 1271 181
rect 1255 147 1345 164
rect 945 100 1345 147
rect -1345 -147 -945 -100
rect -1345 -164 -1255 -147
rect -1271 -181 -1255 -164
rect -1035 -164 -945 -147
rect -887 -147 -487 -100
rect -887 -164 -797 -147
rect -1035 -181 -1019 -164
rect -1271 -197 -1019 -181
rect -813 -181 -797 -164
rect -577 -164 -487 -147
rect -429 -147 -29 -100
rect -429 -164 -339 -147
rect -577 -181 -561 -164
rect -813 -197 -561 -181
rect -355 -181 -339 -164
rect -119 -164 -29 -147
rect 29 -147 429 -100
rect 29 -164 119 -147
rect -119 -181 -103 -164
rect -355 -197 -103 -181
rect 103 -181 119 -164
rect 339 -164 429 -147
rect 487 -147 887 -100
rect 487 -164 577 -147
rect 339 -181 355 -164
rect 103 -197 355 -181
rect 561 -181 577 -164
rect 797 -164 887 -147
rect 945 -147 1345 -100
rect 945 -164 1035 -147
rect 797 -181 813 -164
rect 561 -197 813 -181
rect 1019 -181 1035 -164
rect 1255 -164 1345 -147
rect 1255 -181 1271 -164
rect 1019 -197 1271 -181
<< polycont >>
rect -1255 147 -1035 181
rect -797 147 -577 181
rect -339 147 -119 181
rect 119 147 339 181
rect 577 147 797 181
rect 1035 147 1255 181
rect -1255 -181 -1035 -147
rect -797 -181 -577 -147
rect -339 -181 -119 -147
rect 119 -181 339 -147
rect 577 -181 797 -147
rect 1035 -181 1255 -147
<< locali >>
rect -1271 147 -1255 181
rect -1035 147 -1019 181
rect -813 147 -797 181
rect -577 147 -561 181
rect -355 147 -339 181
rect -119 147 -103 181
rect 103 147 119 181
rect 339 147 355 181
rect 561 147 577 181
rect 797 147 813 181
rect 1019 147 1035 181
rect 1255 147 1271 181
rect -1391 88 -1357 104
rect -1391 -104 -1357 -88
rect -933 88 -899 104
rect -933 -104 -899 -88
rect -475 88 -441 104
rect -475 -104 -441 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 441 88 475 104
rect 441 -104 475 -88
rect 899 88 933 104
rect 899 -104 933 -88
rect 1357 88 1391 104
rect 1357 -104 1391 -88
rect -1271 -181 -1255 -147
rect -1035 -181 -1019 -147
rect -813 -181 -797 -147
rect -577 -181 -561 -147
rect -355 -181 -339 -147
rect -119 -181 -103 -147
rect 103 -181 119 -147
rect 339 -181 355 -147
rect 561 -181 577 -147
rect 797 -181 813 -147
rect 1019 -181 1035 -147
rect 1255 -181 1271 -147
<< viali >>
rect -1237 147 -1053 181
rect -779 147 -595 181
rect -321 147 -137 181
rect 137 147 321 181
rect 595 147 779 181
rect 1053 147 1237 181
rect -1391 -88 -1357 88
rect -933 -88 -899 88
rect -475 -88 -441 88
rect -17 -88 17 88
rect 441 -88 475 88
rect 899 -88 933 88
rect 1357 -88 1391 88
rect -1237 -181 -1053 -147
rect -779 -181 -595 -147
rect -321 -181 -137 -147
rect 137 -181 321 -147
rect 595 -181 779 -147
rect 1053 -181 1237 -147
<< metal1 >>
rect -1249 181 -1041 187
rect -1249 147 -1237 181
rect -1053 147 -1041 181
rect -1249 141 -1041 147
rect -791 181 -583 187
rect -791 147 -779 181
rect -595 147 -583 181
rect -791 141 -583 147
rect -333 181 -125 187
rect -333 147 -321 181
rect -137 147 -125 181
rect -333 141 -125 147
rect 125 181 333 187
rect 125 147 137 181
rect 321 147 333 181
rect 125 141 333 147
rect 583 181 791 187
rect 583 147 595 181
rect 779 147 791 181
rect 583 141 791 147
rect 1041 181 1249 187
rect 1041 147 1053 181
rect 1237 147 1249 181
rect 1041 141 1249 147
rect -1397 88 -1351 100
rect -1397 -88 -1391 88
rect -1357 -88 -1351 88
rect -1397 -100 -1351 -88
rect -939 88 -893 100
rect -939 -88 -933 88
rect -899 -88 -893 88
rect -939 -100 -893 -88
rect -481 88 -435 100
rect -481 -88 -475 88
rect -441 -88 -435 88
rect -481 -100 -435 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 435 88 481 100
rect 435 -88 441 88
rect 475 -88 481 88
rect 435 -100 481 -88
rect 893 88 939 100
rect 893 -88 899 88
rect 933 -88 939 88
rect 893 -100 939 -88
rect 1351 88 1397 100
rect 1351 -88 1357 88
rect 1391 -88 1397 88
rect 1351 -100 1397 -88
rect -1249 -147 -1041 -141
rect -1249 -181 -1237 -147
rect -1053 -181 -1041 -147
rect -1249 -187 -1041 -181
rect -791 -147 -583 -141
rect -791 -181 -779 -147
rect -595 -181 -583 -147
rect -791 -187 -583 -181
rect -333 -147 -125 -141
rect -333 -181 -321 -147
rect -137 -181 -125 -147
rect -333 -187 -125 -181
rect 125 -147 333 -141
rect 125 -181 137 -147
rect 321 -181 333 -147
rect 125 -187 333 -181
rect 583 -147 791 -141
rect 583 -181 595 -147
rect 779 -181 791 -147
rect 583 -187 791 -181
rect 1041 -147 1249 -141
rect 1041 -181 1053 -147
rect 1237 -181 1249 -147
rect 1041 -187 1249 -181
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 1 l 2 m 1 nf 6 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>

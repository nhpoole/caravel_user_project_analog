magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nwell >>
rect 15390 -1694 24486 2310
rect 25972 1912 31856 2230
rect 25972 -1694 32316 1912
<< pwell >>
rect 15390 2474 24486 4420
rect 31466 4346 32270 4350
rect 25972 2400 32270 4346
rect 25972 2394 32268 2400
rect 31460 2286 32268 2394
<< psubdiff >>
rect 15426 4210 15588 4310
rect 24288 4210 24450 4310
rect 15426 4148 15526 4210
rect 15426 2610 15526 2672
rect 24350 4148 24450 4210
rect 24350 2610 24450 2672
rect 15426 2510 15588 2610
rect 24288 2510 24450 2610
rect 26008 4210 26170 4310
rect 31290 4210 31452 4310
rect 26008 4148 26108 4210
rect 26008 2530 26108 2592
rect 31352 4148 31452 4210
rect 31352 2530 31452 2592
rect 26008 2430 26170 2530
rect 31290 2430 31452 2530
<< nsubdiff >>
rect 15426 2174 15588 2274
rect 24288 2174 24450 2274
rect 15426 2112 15526 2174
rect 15426 -1558 15526 -1496
rect 24350 2112 24450 2174
rect 24350 -1558 24450 -1496
rect 15426 -1658 15588 -1558
rect 24288 -1658 24450 -1558
rect 26008 2094 26170 2194
rect 31290 2094 31452 2194
rect 26008 2032 26108 2094
rect 26008 -1558 26108 -1496
rect 31352 2032 31452 2094
rect 31352 -1558 31452 -1496
rect 26008 -1658 26170 -1558
rect 31290 -1658 31452 -1558
<< psubdiffcont >>
rect 15588 4210 24288 4310
rect 15426 2672 15526 4148
rect 24350 2672 24450 4148
rect 15588 2510 24288 2610
rect 26170 4210 31290 4310
rect 26008 2592 26108 4148
rect 31352 2592 31452 4148
rect 26170 2430 31290 2530
<< nsubdiffcont >>
rect 15588 2174 24288 2274
rect 15426 -1496 15526 2112
rect 24350 -1496 24450 2112
rect 15588 -1658 24288 -1558
rect 26170 2094 31290 2194
rect 26008 -1496 26108 2032
rect 31352 -1496 31452 2032
rect 26170 -1658 31290 -1558
<< locali >>
rect 15426 4148 15526 4310
rect 15426 2510 15526 2672
rect 24350 4148 24450 4310
rect 24350 2510 24450 2672
rect 26008 4148 26108 4310
rect 26008 2430 26108 2592
rect 31352 4148 31452 4310
rect 31352 2430 31452 2592
rect 15426 2112 15526 2274
rect 15426 -1658 15526 -1496
rect 24350 2112 24450 2274
rect 24350 -1658 24450 -1496
rect 26008 2032 26108 2194
rect 26008 -1658 26108 -1496
rect 31352 2032 31452 2194
rect 31352 -1658 31452 -1496
<< viali >>
rect 15526 4210 15588 4310
rect 15588 4210 24288 4310
rect 24288 4210 24350 4310
rect 15426 2698 15526 4122
rect 24350 2698 24450 4122
rect 15526 2510 15588 2610
rect 15588 2510 24288 2610
rect 24288 2510 24350 2610
rect 26108 4210 26170 4310
rect 26170 4210 31290 4310
rect 31290 4210 31352 4310
rect 26008 2614 26108 4126
rect 31352 2614 31452 4126
rect 26108 2430 26170 2530
rect 26170 2430 31290 2530
rect 31290 2430 31352 2530
rect 15526 2174 15588 2274
rect 15588 2174 24288 2274
rect 24288 2174 24350 2274
rect 15426 -1360 15526 1976
rect 31606 2226 31654 2274
rect 31712 2228 31760 2276
rect 31848 2228 31896 2276
rect 32204 2228 32252 2276
rect 24350 -1360 24450 1976
rect 15526 -1658 15588 -1558
rect 15588 -1658 24288 -1558
rect 24288 -1658 24350 -1558
rect 26108 2094 26170 2194
rect 26170 2094 31290 2194
rect 31290 2094 31352 2194
rect 26008 -1375 26108 1911
rect 31352 -1375 31452 1911
rect 26108 -1658 26170 -1558
rect 26170 -1658 31290 -1558
rect 31290 -1658 31352 -1558
<< metal1 >>
rect 15420 4310 24456 4316
rect 15420 4210 15526 4310
rect 24350 4210 24456 4310
rect 15420 4204 24456 4210
rect 15420 4122 15532 4204
rect 15420 2698 15426 4122
rect 15526 2698 15532 4122
rect 15914 3904 15924 4204
rect 23656 3904 23666 4204
rect 24344 4122 24456 4204
rect 17550 3726 22522 3756
rect 17550 3640 17600 3726
rect 17696 3640 18180 3726
rect 18276 3640 18780 3726
rect 18876 3640 19380 3726
rect 19476 3640 19980 3726
rect 20076 3640 20580 3726
rect 20676 3640 21180 3726
rect 21276 3640 21780 3726
rect 21876 3640 22380 3726
rect 22476 3640 22522 3726
rect 17550 3612 22522 3640
rect 17614 3202 17674 3612
rect 17854 3282 17914 3612
rect 18304 3388 21514 3448
rect 21574 3388 21580 3448
rect 18304 3282 18364 3388
rect 18766 3292 18826 3388
rect 19220 3286 19280 3388
rect 19682 3286 19742 3388
rect 20136 3286 20196 3388
rect 20586 3292 20646 3388
rect 21052 3298 21112 3388
rect 21508 3292 21568 3388
rect 21742 3204 21802 3612
rect 21968 3280 22028 3612
rect 15420 2616 15532 2698
rect 17622 2616 17682 3076
rect 17850 2616 17910 3006
rect 18078 2768 18138 3084
rect 18310 2894 18376 3006
rect 18772 2894 18838 3006
rect 19226 2894 19292 3006
rect 19688 2894 19754 3006
rect 20142 2894 20208 3006
rect 20592 2894 20658 3006
rect 21058 2894 21124 3006
rect 21514 2894 21580 3006
rect 18310 2828 21580 2894
rect 18078 2702 18138 2708
rect 21748 2616 21808 3076
rect 21976 2616 22036 3008
rect 22208 2616 22268 3612
rect 24344 2698 24350 4122
rect 24450 2698 24456 4122
rect 24344 2616 24456 2698
rect 15420 2610 24456 2616
rect 15420 2510 15526 2610
rect 24350 2510 24456 2610
rect 15420 2504 24456 2510
rect 26002 4310 31458 4316
rect 26002 4210 26108 4310
rect 31352 4210 31458 4310
rect 26002 4204 31458 4210
rect 26002 4126 26114 4204
rect 26002 2614 26008 4126
rect 26108 2614 26114 4126
rect 26714 3904 26724 4204
rect 30736 3904 30746 4204
rect 31346 4126 31458 4204
rect 26312 3726 31284 3756
rect 26312 3640 26362 3726
rect 26458 3640 26942 3726
rect 27038 3640 27542 3726
rect 27638 3640 28142 3726
rect 28238 3640 28742 3726
rect 28838 3640 29342 3726
rect 29438 3640 29942 3726
rect 30038 3640 30542 3726
rect 30638 3640 31142 3726
rect 31238 3640 31284 3726
rect 26312 3612 31284 3640
rect 26376 3202 26436 3612
rect 26616 3282 26676 3612
rect 26002 2536 26114 2614
rect 26384 2536 26444 3076
rect 26612 2536 26672 3006
rect 26840 2536 26900 3612
rect 27066 3388 30330 3448
rect 27066 3282 27126 3388
rect 27528 3292 27588 3388
rect 27982 3286 28042 3388
rect 28444 3286 28504 3388
rect 28898 3286 28958 3388
rect 29348 3292 29408 3388
rect 29814 3298 29874 3388
rect 30270 3292 30330 3388
rect 30730 3280 30790 3612
rect 27066 2894 27126 3002
rect 27528 2894 27588 3004
rect 27982 2896 28042 3004
rect 27976 2894 27982 2896
rect 27059 2834 27066 2894
rect 27126 2834 27528 2894
rect 27588 2836 27982 2894
rect 28042 2894 28048 2896
rect 28444 2894 28504 3006
rect 28898 2894 28958 3006
rect 29348 2894 29408 3006
rect 29814 2894 29874 3002
rect 30270 2894 30330 3006
rect 28042 2836 28444 2894
rect 27588 2834 28444 2836
rect 28504 2834 28898 2894
rect 28958 2834 29348 2894
rect 29408 2834 29814 2894
rect 29874 2834 30270 2894
rect 30330 2834 30337 2894
rect 27059 2828 30337 2834
rect 30504 2686 30564 3110
rect 30498 2626 30504 2686
rect 30564 2626 30570 2686
rect 30738 2536 30798 3008
rect 30970 2536 31030 3612
rect 31346 2614 31352 4126
rect 31452 2614 31458 4126
rect 31346 2538 31458 2614
rect 31346 2536 31542 2538
rect 26002 2530 31542 2536
rect 26002 2430 26108 2530
rect 31352 2442 31542 2530
rect 31352 2430 31458 2442
rect 26002 2424 31458 2430
rect 30504 2344 30564 2350
rect 25234 2284 30504 2344
rect 30564 2284 31566 2344
rect 15420 2274 24456 2280
rect 15420 2174 15526 2274
rect 24350 2174 24456 2274
rect 15420 2168 24456 2174
rect 15420 1976 15532 2168
rect 15420 -1360 15426 1976
rect 15526 1614 15532 1976
rect 15790 1614 15850 2168
rect 16018 1614 16078 2168
rect 16244 1614 16304 2168
rect 16702 2026 23178 2086
rect 15526 1554 16304 1614
rect 16468 1554 16474 1614
rect 16534 1554 16540 1614
rect 15526 -1360 15532 1554
rect 15790 1322 15850 1554
rect 16018 1438 16078 1554
rect 16244 1338 16304 1554
rect 16474 1446 16534 1554
rect 16702 1298 16762 2026
rect 17620 1902 22264 1962
rect 16924 1554 16930 1614
rect 16990 1554 16996 1614
rect 17384 1554 17390 1614
rect 17450 1554 17456 1614
rect 16930 1448 16990 1554
rect 17390 1442 17450 1554
rect 17620 1304 17680 1902
rect 18528 1778 21344 1838
rect 17840 1554 17846 1614
rect 17906 1554 17912 1614
rect 18298 1554 18304 1614
rect 18364 1554 18370 1614
rect 17846 1448 17906 1554
rect 18304 1448 18364 1554
rect 18528 1310 18588 1778
rect 19452 1662 20430 1722
rect 18762 1554 18768 1614
rect 18828 1554 18834 1614
rect 19216 1554 19222 1614
rect 19282 1554 19288 1614
rect 18768 1444 18828 1554
rect 19222 1442 19282 1554
rect 19452 1302 19512 1662
rect 19676 1554 19682 1614
rect 19742 1554 19748 1614
rect 19906 1554 19912 1614
rect 19972 1554 19978 1614
rect 20134 1554 20140 1614
rect 20200 1554 20206 1614
rect 19682 1444 19742 1554
rect 19912 1332 19972 1554
rect 20140 1436 20200 1554
rect 20370 1354 20430 1662
rect 20590 1554 20596 1614
rect 20656 1554 20662 1614
rect 21050 1554 21056 1614
rect 21116 1554 21122 1614
rect 20596 1442 20656 1554
rect 21056 1448 21116 1554
rect 21284 1350 21344 1778
rect 21506 1554 21512 1614
rect 21572 1554 21578 1614
rect 21962 1554 21968 1614
rect 22028 1554 22034 1614
rect 21512 1448 21572 1554
rect 21968 1448 22028 1554
rect 22204 1314 22264 1902
rect 22418 1554 22424 1614
rect 22484 1554 22490 1614
rect 22876 1554 22882 1614
rect 22942 1554 22948 1614
rect 22424 1452 22484 1554
rect 22882 1448 22942 1554
rect 23118 1322 23178 2026
rect 23572 1614 23632 2168
rect 23804 1614 23864 2168
rect 24030 1614 24090 2168
rect 24344 1976 24456 2168
rect 24344 1614 24350 1976
rect 23336 1554 23342 1614
rect 23402 1554 23408 1614
rect 23572 1554 24350 1614
rect 23342 1444 23402 1554
rect 23572 1320 23632 1554
rect 23804 1440 23864 1554
rect 24030 1338 24090 1554
rect 15788 -982 15848 -162
rect 16020 -982 16080 -254
rect 16246 -982 16306 -130
rect 16478 -360 16538 -252
rect 16934 -360 16994 -254
rect 16472 -420 16478 -360
rect 16538 -420 16544 -360
rect 16928 -420 16934 -360
rect 16994 -420 17000 -360
rect 17162 -728 17222 -136
rect 17394 -360 17454 -248
rect 17850 -360 17910 -254
rect 17388 -420 17394 -360
rect 17454 -420 17460 -360
rect 17844 -420 17850 -360
rect 17910 -420 17916 -360
rect 18078 -594 18138 -134
rect 18308 -360 18368 -254
rect 18772 -360 18832 -250
rect 18302 -420 18308 -360
rect 18368 -420 18374 -360
rect 18766 -420 18772 -360
rect 18832 -420 18838 -360
rect 18994 -470 19054 -116
rect 19222 -360 19282 -256
rect 19678 -360 19738 -256
rect 20146 -360 20206 -256
rect 20604 -360 20664 -260
rect 19216 -420 19222 -360
rect 19282 -420 19288 -360
rect 19672 -420 19678 -360
rect 19738 -420 19744 -360
rect 20140 -420 20146 -360
rect 20206 -420 20212 -360
rect 20598 -420 20604 -360
rect 20664 -420 20670 -360
rect 20824 -470 20884 -150
rect 21060 -360 21120 -254
rect 21516 -360 21576 -254
rect 21054 -420 21060 -360
rect 21120 -420 21126 -360
rect 21510 -420 21516 -360
rect 21576 -420 21582 -360
rect 18994 -530 20884 -470
rect 21740 -594 21800 -136
rect 21972 -360 22032 -254
rect 22428 -360 22488 -258
rect 21966 -420 21972 -360
rect 22032 -420 22038 -360
rect 22422 -420 22428 -360
rect 22488 -420 22494 -360
rect 18078 -654 21800 -594
rect 22660 -728 22720 -138
rect 22886 -360 22946 -254
rect 23346 -360 23406 -250
rect 22880 -420 22886 -360
rect 22946 -420 22952 -360
rect 23340 -420 23346 -360
rect 23406 -420 23412 -360
rect 17162 -788 22720 -728
rect 23576 -982 23636 -118
rect 23806 -982 23866 -252
rect 24034 -982 24094 -124
rect 24344 -982 24350 1554
rect 15760 -992 24350 -982
rect 15760 -1078 15774 -992
rect 15870 -1078 16374 -992
rect 16470 -1078 16974 -992
rect 17070 -1078 17574 -992
rect 17670 -1078 18174 -992
rect 18270 -1078 18774 -992
rect 18870 -1078 19374 -992
rect 19470 -1078 19974 -992
rect 20070 -1078 20574 -992
rect 20670 -1078 21174 -992
rect 21270 -1078 21774 -992
rect 21870 -1078 22374 -992
rect 22470 -1078 22974 -992
rect 23070 -1078 23574 -992
rect 23670 -1078 23994 -992
rect 24090 -1078 24350 -992
rect 15760 -1092 24350 -1078
rect 15420 -1552 15532 -1360
rect 15914 -1552 15924 -1252
rect 23656 -1552 23666 -1252
rect 24344 -1360 24350 -1092
rect 24450 -982 24456 1976
rect 24450 -1092 24458 -982
rect 24450 -1360 24456 -1092
rect 24344 -1552 24456 -1360
rect 15420 -1558 24456 -1552
rect 15420 -1658 15526 -1558
rect 24350 -1658 24456 -1558
rect 15420 -1664 24456 -1658
rect 25234 -5664 25294 2284
rect 30504 2278 30564 2284
rect 31506 2280 31566 2284
rect 31506 2274 31666 2280
rect 31506 2226 31606 2274
rect 31654 2226 31666 2274
rect 31506 2220 31666 2226
rect 31700 2276 31908 2282
rect 31700 2228 31712 2276
rect 31760 2228 31848 2276
rect 31896 2228 31908 2276
rect 31700 2222 31908 2228
rect 32192 2276 32478 2282
rect 32192 2228 32204 2276
rect 32252 2228 32478 2276
rect 32192 2222 32478 2228
rect 25546 2200 25606 2206
rect 25400 -420 25406 -360
rect 25466 -420 25472 -360
rect 25406 -3260 25466 -420
rect 25406 -3266 25468 -3260
rect 25406 -3326 25408 -3266
rect 25406 -3332 25468 -3326
rect 25228 -5724 25234 -5664
rect 25294 -5724 25300 -5664
rect 15000 -5988 15124 -5928
rect 15184 -5988 15190 -5928
rect 15010 -9710 15116 -9650
rect 15176 -9710 15182 -9650
rect 23994 -11954 24062 -11894
rect 24122 -11954 24128 -11894
rect 25406 -16304 25466 -3332
rect 25546 -9650 25606 2140
rect 26002 2194 31458 2200
rect 26002 2094 26108 2194
rect 31352 2094 31458 2194
rect 26002 2088 31458 2094
rect 26002 1911 26114 2088
rect 26002 -982 26008 1911
rect 26000 -1092 26008 -982
rect 26002 -1375 26008 -1092
rect 26108 420 26114 1911
rect 26384 1778 26444 2088
rect 26612 1858 26672 2088
rect 26384 420 26444 670
rect 26612 420 26672 562
rect 26842 420 26902 2088
rect 30504 2032 30564 2038
rect 27066 2026 27126 2032
rect 27528 2026 27588 2032
rect 27982 2026 28042 2032
rect 28444 2026 28504 2032
rect 28898 2026 28958 2032
rect 29348 2026 29408 2032
rect 29814 2026 29874 2032
rect 30270 2026 30330 2032
rect 27060 1966 27066 2026
rect 27126 1966 27528 2026
rect 27588 1966 27982 2026
rect 28042 1966 28444 2026
rect 28504 1966 28898 2026
rect 28958 1966 29348 2026
rect 29408 1966 29814 2026
rect 29874 1966 30270 2026
rect 30330 1966 30336 2026
rect 27066 1854 27126 1966
rect 27528 1870 27588 1966
rect 27982 1864 28042 1966
rect 28444 1864 28504 1966
rect 28898 1864 28958 1966
rect 29348 1870 29408 1966
rect 29814 1876 29874 1966
rect 30270 1870 30330 1966
rect 30504 1732 30564 1972
rect 30734 1856 30794 2088
rect 30962 1764 31022 2088
rect 31346 1994 31458 2088
rect 31346 1911 31542 1994
rect 26108 360 26902 420
rect 27074 454 27134 566
rect 27536 454 27596 550
rect 27990 454 28050 556
rect 28452 454 28512 556
rect 28906 454 28966 556
rect 29356 454 29416 550
rect 29822 454 29882 544
rect 30278 454 30338 550
rect 30734 472 30794 562
rect 30964 472 31024 638
rect 31346 472 31352 1911
rect 27074 394 30278 454
rect 30338 394 30344 454
rect 30734 412 31352 472
rect 26108 -982 26114 360
rect 26384 -982 26444 360
rect 26612 -982 26672 360
rect 26842 -982 26902 360
rect 30734 -982 30794 412
rect 30964 -982 31024 412
rect 26108 -992 31274 -982
rect 26108 -1078 26290 -992
rect 26386 -1078 26890 -992
rect 26986 -1078 27490 -992
rect 27586 -1078 28090 -992
rect 28186 -1078 28690 -992
rect 28786 -1078 29290 -992
rect 29386 -1078 29890 -992
rect 29986 -1078 30490 -992
rect 30586 -1078 31090 -992
rect 31186 -1078 31274 -992
rect 26108 -1092 31274 -1078
rect 26108 -1375 26114 -1092
rect 26002 -1552 26114 -1375
rect 26714 -1552 26724 -1252
rect 30736 -1552 30746 -1252
rect 31346 -1375 31352 412
rect 31452 1898 31542 1911
rect 31452 -1375 31458 1898
rect 31346 -1552 31458 -1375
rect 26002 -1558 31458 -1552
rect 26002 -1658 26108 -1558
rect 31352 -1658 31458 -1558
rect 26002 -1664 31458 -1658
rect 26914 -9650 26974 -9644
rect 25540 -9710 25546 -9650
rect 25606 -9710 25612 -9650
rect 25406 -23240 25466 -16364
rect 25546 -11894 25606 -9710
rect 26914 -9716 26974 -9710
rect 25400 -23300 25406 -23240
rect 25466 -23300 25472 -23240
rect 15118 -27650 15178 -27644
rect 25546 -27650 25606 -11954
rect 35856 -11894 35916 -11888
rect 35916 -11954 36076 -11894
rect 35856 -11960 35916 -11954
rect 25540 -27710 25546 -27650
rect 25606 -27710 25612 -27650
rect 26908 -27710 26914 -27650
rect 26974 -27710 27050 -27650
rect 15118 -27716 15178 -27710
<< via1 >>
rect 15532 3904 15914 4204
rect 23666 3904 24344 4204
rect 17600 3640 17696 3726
rect 18180 3640 18276 3726
rect 18780 3640 18876 3726
rect 19380 3640 19476 3726
rect 19980 3640 20076 3726
rect 20580 3640 20676 3726
rect 21180 3640 21276 3726
rect 21780 3640 21876 3726
rect 22380 3640 22476 3726
rect 21514 3388 21574 3448
rect 18078 2708 18138 2768
rect 26114 3904 26714 4204
rect 30746 3904 31346 4204
rect 26362 3640 26458 3726
rect 26942 3640 27038 3726
rect 27542 3640 27638 3726
rect 28142 3640 28238 3726
rect 28742 3640 28838 3726
rect 29342 3640 29438 3726
rect 29942 3640 30038 3726
rect 30542 3640 30638 3726
rect 31142 3640 31238 3726
rect 27066 2834 27126 2894
rect 27528 2834 27588 2894
rect 27982 2836 28042 2896
rect 28444 2834 28504 2894
rect 28898 2834 28958 2894
rect 29348 2834 29408 2894
rect 29814 2834 29874 2894
rect 30270 2834 30330 2894
rect 30504 2626 30564 2686
rect 30504 2284 30564 2344
rect 16474 1554 16534 1614
rect 16930 1554 16990 1614
rect 17390 1554 17450 1614
rect 17846 1554 17906 1614
rect 18304 1554 18364 1614
rect 18768 1554 18828 1614
rect 19222 1554 19282 1614
rect 19682 1554 19742 1614
rect 19912 1554 19972 1614
rect 20140 1554 20200 1614
rect 20596 1554 20656 1614
rect 21056 1554 21116 1614
rect 21512 1554 21572 1614
rect 21968 1554 22028 1614
rect 22424 1554 22484 1614
rect 22882 1554 22942 1614
rect 23342 1554 23402 1614
rect 16478 -420 16538 -360
rect 16934 -420 16994 -360
rect 17394 -420 17454 -360
rect 17850 -420 17910 -360
rect 18308 -420 18368 -360
rect 18772 -420 18832 -360
rect 19222 -420 19282 -360
rect 19678 -420 19738 -360
rect 20146 -420 20206 -360
rect 20604 -420 20664 -360
rect 21060 -420 21120 -360
rect 21516 -420 21576 -360
rect 21972 -420 22032 -360
rect 22428 -420 22488 -360
rect 22886 -420 22946 -360
rect 23346 -420 23406 -360
rect 15774 -1078 15870 -992
rect 16374 -1078 16470 -992
rect 16974 -1078 17070 -992
rect 17574 -1078 17670 -992
rect 18174 -1078 18270 -992
rect 18774 -1078 18870 -992
rect 19374 -1078 19470 -992
rect 19974 -1078 20070 -992
rect 20574 -1078 20670 -992
rect 21174 -1078 21270 -992
rect 21774 -1078 21870 -992
rect 22374 -1078 22470 -992
rect 22974 -1078 23070 -992
rect 23574 -1078 23670 -992
rect 23994 -1078 24090 -992
rect 15532 -1552 15914 -1252
rect 23666 -1552 24344 -1252
rect 25546 2140 25606 2200
rect 25406 -420 25466 -360
rect 25408 -3326 25468 -3266
rect 25234 -5724 25294 -5664
rect 15124 -5988 15184 -5928
rect 15116 -9710 15176 -9650
rect 24062 -11954 24122 -11894
rect 27066 1966 27126 2026
rect 27528 1966 27588 2026
rect 27982 1966 28042 2026
rect 28444 1966 28504 2026
rect 28898 1966 28958 2026
rect 29348 1966 29408 2026
rect 29814 1966 29874 2026
rect 30270 1966 30330 2026
rect 30504 1972 30564 2032
rect 30278 394 30338 454
rect 26290 -1078 26386 -992
rect 26890 -1078 26986 -992
rect 27490 -1078 27586 -992
rect 28090 -1078 28186 -992
rect 28690 -1078 28786 -992
rect 29290 -1078 29386 -992
rect 29890 -1078 29986 -992
rect 30490 -1078 30586 -992
rect 31090 -1078 31186 -992
rect 26114 -1552 26714 -1252
rect 30746 -1552 31346 -1252
rect 25546 -9710 25606 -9650
rect 26914 -9710 26974 -9650
rect 25406 -16364 25466 -16304
rect 25546 -11954 25606 -11894
rect 25406 -23300 25466 -23240
rect 35856 -11954 35916 -11894
rect 15118 -27710 15178 -27650
rect 25546 -27710 25606 -27650
rect 26914 -27710 26974 -27650
<< metal2 >>
rect 15532 4204 15914 4214
rect 15532 3894 15914 3904
rect 23666 4204 24344 4214
rect 23666 3894 24344 3904
rect 26114 4204 26714 4214
rect 26114 3894 26714 3904
rect 30746 4204 31346 4214
rect 30746 3894 31346 3904
rect 17550 3726 22522 3756
rect 17550 3640 17600 3726
rect 17696 3640 18180 3726
rect 18276 3640 18780 3726
rect 18876 3640 19380 3726
rect 19476 3640 19980 3726
rect 20076 3640 20580 3726
rect 20676 3640 21180 3726
rect 21276 3640 21780 3726
rect 21876 3640 22380 3726
rect 22476 3640 22522 3726
rect 17550 3612 22522 3640
rect 26312 3726 31284 3756
rect 26312 3640 26362 3726
rect 26458 3640 26942 3726
rect 27038 3640 27542 3726
rect 27638 3640 28142 3726
rect 28238 3640 28742 3726
rect 28838 3640 29342 3726
rect 29438 3640 29942 3726
rect 30038 3640 30542 3726
rect 30638 3640 31142 3726
rect 31238 3640 31284 3726
rect 26312 3612 31284 3640
rect 21514 3448 21574 3454
rect 21574 3388 25606 3448
rect 21514 3382 21574 3388
rect 18072 2708 18078 2768
rect 18138 2708 18144 2768
rect 16474 1614 16534 1620
rect 16930 1614 16990 1620
rect 17390 1614 17450 1620
rect 17846 1614 17906 1620
rect 18078 1614 18138 2708
rect 25546 2200 25606 3388
rect 27066 2894 27126 2900
rect 25540 2140 25546 2200
rect 25606 2140 25612 2200
rect 27066 2026 27126 2834
rect 27066 1960 27126 1966
rect 27528 2894 27588 2900
rect 27528 2026 27588 2834
rect 27982 2896 28042 2902
rect 27982 2026 28042 2836
rect 28444 2894 28504 2900
rect 28444 2026 28504 2834
rect 28898 2894 28958 2900
rect 28898 2026 28958 2834
rect 29348 2894 29408 2900
rect 29348 2026 29408 2834
rect 29814 2894 29874 2900
rect 29814 2026 29874 2834
rect 30270 2894 30330 2900
rect 30270 2026 30330 2834
rect 30504 2686 30564 2692
rect 30504 2344 30564 2626
rect 30498 2284 30504 2344
rect 30564 2284 30570 2344
rect 30504 2032 30564 2284
rect 27976 1966 27982 2026
rect 28042 1966 28048 2026
rect 28438 1966 28444 2026
rect 28504 1966 28510 2026
rect 29342 1966 29348 2026
rect 29408 1966 29414 2026
rect 29808 1966 29814 2026
rect 29874 1966 29880 2026
rect 30498 1972 30504 2032
rect 30564 1972 30570 2032
rect 27528 1960 27588 1966
rect 28898 1960 28958 1966
rect 30270 1960 30330 1966
rect 18304 1614 18364 1620
rect 18768 1614 18828 1620
rect 19222 1614 19282 1620
rect 19682 1614 19742 1620
rect 19912 1614 19972 1620
rect 20140 1614 20200 1620
rect 20596 1614 20656 1620
rect 21056 1614 21116 1620
rect 21512 1614 21572 1620
rect 21968 1614 22028 1620
rect 22424 1614 22484 1620
rect 22882 1614 22942 1620
rect 23342 1614 23402 1620
rect 16534 1554 16930 1614
rect 16990 1554 17390 1614
rect 17450 1554 17846 1614
rect 17906 1554 18304 1614
rect 18364 1554 18768 1614
rect 18828 1554 19222 1614
rect 19282 1554 19682 1614
rect 19742 1554 19912 1614
rect 19972 1554 20140 1614
rect 20200 1554 20596 1614
rect 20656 1554 21056 1614
rect 21116 1554 21512 1614
rect 21572 1554 21968 1614
rect 22028 1554 22424 1614
rect 22484 1554 22882 1614
rect 22942 1554 23342 1614
rect 16474 1548 16534 1554
rect 16930 1548 16990 1554
rect 17390 1548 17450 1554
rect 17846 1548 17906 1554
rect 18304 1548 18364 1554
rect 18768 1548 18828 1554
rect 19222 1548 19282 1554
rect 19682 1548 19742 1554
rect 19912 1548 19972 1554
rect 20140 1548 20200 1554
rect 20596 1548 20656 1554
rect 21056 1548 21116 1554
rect 21512 1548 21572 1554
rect 21968 1548 22028 1554
rect 22424 1548 22484 1554
rect 22882 1548 22942 1554
rect 23342 1548 23402 1554
rect 30278 454 30338 460
rect 30338 394 31902 454
rect 30278 388 30338 394
rect 16478 -360 16538 -354
rect 16934 -360 16994 -354
rect 17394 -360 17454 -354
rect 17850 -360 17910 -354
rect 18308 -360 18368 -354
rect 18772 -360 18832 -354
rect 19222 -360 19282 -354
rect 19678 -360 19738 -354
rect 20146 -360 20206 -354
rect 20604 -360 20664 -354
rect 21060 -360 21120 -354
rect 21516 -360 21576 -354
rect 21972 -360 22032 -354
rect 22428 -360 22488 -354
rect 22886 -360 22946 -354
rect 23346 -360 23406 -354
rect 25406 -360 25466 -354
rect 16538 -420 16934 -360
rect 16994 -420 17394 -360
rect 17454 -420 17850 -360
rect 17910 -420 18308 -360
rect 18368 -420 18772 -360
rect 18832 -420 19222 -360
rect 19282 -420 19678 -360
rect 19738 -420 20146 -360
rect 20206 -420 20604 -360
rect 20664 -420 21060 -360
rect 21120 -420 21516 -360
rect 21576 -420 21972 -360
rect 22032 -420 22428 -360
rect 22488 -420 22886 -360
rect 22946 -420 23346 -360
rect 23406 -420 25406 -360
rect 16478 -426 16538 -420
rect 16934 -426 16994 -420
rect 17394 -426 17454 -420
rect 17850 -426 17910 -420
rect 18308 -426 18368 -420
rect 18772 -426 18832 -420
rect 19222 -426 19282 -420
rect 19678 -426 19738 -420
rect 20146 -426 20206 -420
rect 20604 -426 20664 -420
rect 21060 -426 21120 -420
rect 21516 -426 21576 -420
rect 21972 -426 22032 -420
rect 22428 -426 22488 -420
rect 22886 -426 22946 -420
rect 23346 -426 23406 -420
rect 25406 -426 25466 -420
rect 31802 -948 31902 394
rect 15760 -992 24116 -982
rect 15760 -1078 15774 -992
rect 15870 -1078 16374 -992
rect 16470 -1078 16974 -992
rect 17070 -1078 17574 -992
rect 17670 -1078 18174 -992
rect 18270 -1078 18774 -992
rect 18870 -1078 19374 -992
rect 19470 -1078 19974 -992
rect 20070 -1078 20574 -992
rect 20670 -1078 21174 -992
rect 21270 -1078 21774 -992
rect 21870 -1078 22374 -992
rect 22470 -1078 22974 -992
rect 23070 -1078 23574 -992
rect 23670 -1078 23994 -992
rect 24090 -1078 24116 -992
rect 15760 -1092 24116 -1078
rect 26276 -992 31274 -982
rect 26276 -1078 26290 -992
rect 26386 -1078 26890 -992
rect 26986 -1078 27490 -992
rect 27586 -1078 28090 -992
rect 28186 -1078 28690 -992
rect 28786 -1078 29290 -992
rect 29386 -1078 29890 -992
rect 29986 -1078 30490 -992
rect 30586 -1078 31090 -992
rect 31186 -1078 31274 -992
rect 31802 -1048 36438 -948
rect 26276 -1092 31274 -1078
rect 15532 -1252 15914 -1242
rect 15532 -1562 15914 -1552
rect 23666 -1252 24344 -1242
rect 23666 -1562 24344 -1552
rect 26114 -1252 26714 -1242
rect 26114 -1562 26714 -1552
rect 30746 -1252 31346 -1242
rect 30746 -1562 31346 -1552
rect 19242 -3326 25408 -3266
rect 25468 -3326 27720 -3266
rect 25234 -5664 25294 -5658
rect 16180 -5724 25234 -5664
rect 15124 -5928 15184 -5922
rect 16180 -5928 16240 -5724
rect 25234 -5730 25294 -5724
rect 15184 -5988 16240 -5928
rect 15124 -5994 15184 -5988
rect 25616 -7958 25676 -7949
rect 25676 -8018 27308 -7958
rect 25616 -8027 25676 -8018
rect 36338 -8128 36438 -1048
rect 15116 -9650 15176 -9644
rect 25546 -9650 25606 -9644
rect 15176 -9710 25546 -9650
rect 25606 -9710 26914 -9650
rect 26974 -9710 26980 -9650
rect 15116 -9716 15176 -9710
rect 25546 -9716 25606 -9710
rect 24062 -11894 24122 -11888
rect 24122 -11954 25546 -11894
rect 25606 -11954 35856 -11894
rect 35916 -11954 35922 -11894
rect 24062 -11960 24122 -11954
rect 10630 -13357 10690 -13352
rect 10600 -13447 10609 -13357
rect 10699 -13447 10708 -13357
rect 10630 -25958 10690 -13447
rect 25300 -13586 25360 -13577
rect 23754 -13646 25300 -13586
rect 38988 -13646 40380 -13586
rect 25300 -13655 25360 -13646
rect 23180 -16364 25406 -16304
rect 25466 -16364 32052 -16304
rect 25406 -23240 25466 -23234
rect 19246 -23300 25406 -23240
rect 25466 -23300 27852 -23240
rect 25406 -23306 25466 -23300
rect 10630 -26018 12078 -25958
rect 25420 -26018 27060 -25958
rect 25420 -26157 25480 -26018
rect 40320 -26157 40380 -13646
rect 25398 -26247 25407 -26157
rect 25497 -26247 25506 -26157
rect 40296 -26247 40305 -26157
rect 40395 -26247 40404 -26157
rect 25420 -26252 25480 -26247
rect 40320 -26252 40380 -26247
rect 25546 -27650 25606 -27644
rect 26914 -27650 26974 -27644
rect 15112 -27710 15118 -27650
rect 15178 -27710 25546 -27650
rect 25606 -27710 26914 -27650
rect 25546 -27716 25606 -27710
rect 26914 -27716 26974 -27710
<< via2 >>
rect 15532 3904 15914 4204
rect 23666 3904 24344 4204
rect 26114 3904 26714 4204
rect 30746 3904 31346 4204
rect 17600 3640 17696 3726
rect 18180 3640 18276 3726
rect 18780 3640 18876 3726
rect 19380 3640 19476 3726
rect 19980 3640 20076 3726
rect 20580 3640 20676 3726
rect 21180 3640 21276 3726
rect 21780 3640 21876 3726
rect 22380 3640 22476 3726
rect 26362 3640 26458 3726
rect 26942 3640 27038 3726
rect 27542 3640 27638 3726
rect 28142 3640 28238 3726
rect 28742 3640 28838 3726
rect 29342 3640 29438 3726
rect 29942 3640 30038 3726
rect 30542 3640 30638 3726
rect 31142 3640 31238 3726
rect 15774 -1078 15870 -992
rect 16374 -1078 16470 -992
rect 16974 -1078 17070 -992
rect 17574 -1078 17670 -992
rect 18174 -1078 18270 -992
rect 18774 -1078 18870 -992
rect 19374 -1078 19470 -992
rect 19974 -1078 20070 -992
rect 20574 -1078 20670 -992
rect 21174 -1078 21270 -992
rect 21774 -1078 21870 -992
rect 22374 -1078 22470 -992
rect 22974 -1078 23070 -992
rect 23574 -1078 23670 -992
rect 23994 -1078 24090 -992
rect 26290 -1078 26386 -992
rect 26890 -1078 26986 -992
rect 27490 -1078 27586 -992
rect 28090 -1078 28186 -992
rect 28690 -1078 28786 -992
rect 29290 -1078 29386 -992
rect 29890 -1078 29986 -992
rect 30490 -1078 30586 -992
rect 31090 -1078 31186 -992
rect 15532 -1552 15914 -1252
rect 23666 -1552 24344 -1252
rect 26114 -1552 26714 -1252
rect 30746 -1552 31346 -1252
rect 25616 -8018 25676 -7958
rect 10609 -13447 10699 -13357
rect 25300 -13646 25360 -13586
rect 25407 -26247 25497 -26157
rect 40305 -26247 40395 -26157
<< metal3 >>
rect 15522 4204 15924 4209
rect 15522 3904 15532 4204
rect 15914 3904 15924 4204
rect 15522 3899 15924 3904
rect 23656 4204 24354 4209
rect 23656 3904 23666 4204
rect 24344 3904 24354 4204
rect 23656 3899 24354 3904
rect 26104 4204 26724 4209
rect 26104 3904 26114 4204
rect 26714 3904 26724 4204
rect 26104 3899 26724 3904
rect 30736 4204 31356 4209
rect 30736 3904 30746 4204
rect 31346 3904 31356 4204
rect 30736 3899 31356 3904
rect 17550 3726 22522 3756
rect 17550 3640 17600 3726
rect 17696 3640 18180 3726
rect 18276 3640 18780 3726
rect 18876 3640 19380 3726
rect 19476 3640 19980 3726
rect 20076 3640 20580 3726
rect 20676 3640 21180 3726
rect 21276 3640 21780 3726
rect 21876 3640 22380 3726
rect 22476 3640 22522 3726
rect 17550 3612 22522 3640
rect 26312 3726 31284 3756
rect 26312 3640 26362 3726
rect 26458 3640 26942 3726
rect 27038 3640 27542 3726
rect 27638 3640 28142 3726
rect 28238 3640 28742 3726
rect 28838 3640 29342 3726
rect 29438 3640 29942 3726
rect 30038 3640 30542 3726
rect 30638 3640 31142 3726
rect 31238 3640 31284 3726
rect 26312 3612 31284 3640
rect 15760 -992 24116 -982
rect 15760 -1078 15774 -992
rect 15870 -1078 16374 -992
rect 16470 -1078 16974 -992
rect 17070 -1078 17574 -992
rect 17670 -1078 18174 -992
rect 18270 -1078 18774 -992
rect 18870 -1078 19374 -992
rect 19470 -1078 19974 -992
rect 20070 -1078 20574 -992
rect 20670 -1078 21174 -992
rect 21270 -1078 21774 -992
rect 21870 -1078 22374 -992
rect 22470 -1078 22974 -992
rect 23070 -1078 23574 -992
rect 23670 -1078 23994 -992
rect 24090 -1078 24116 -992
rect 15760 -1092 24116 -1078
rect 26276 -992 31274 -982
rect 26276 -1078 26290 -992
rect 26386 -1078 26890 -992
rect 26986 -1078 27490 -992
rect 27586 -1078 28090 -992
rect 28186 -1078 28690 -992
rect 28786 -1078 29290 -992
rect 29386 -1078 29890 -992
rect 29986 -1078 30490 -992
rect 30586 -1078 31090 -992
rect 31186 -1078 31274 -992
rect 26276 -1092 31274 -1078
rect 15522 -1252 15924 -1247
rect 15522 -1552 15532 -1252
rect 15914 -1552 15924 -1252
rect 15522 -1557 15924 -1552
rect 23656 -1252 24354 -1247
rect 23656 -1552 23666 -1252
rect 24344 -1552 24354 -1252
rect 23656 -1557 24354 -1552
rect 26104 -1252 26724 -1247
rect 26104 -1552 26114 -1252
rect 26714 -1552 26724 -1252
rect 26104 -1557 26724 -1552
rect 30736 -1252 31356 -1247
rect 30736 -1552 30746 -1252
rect 31346 -1552 31356 -1252
rect 30736 -1557 31356 -1552
rect 25611 -7958 25681 -7953
rect 25596 -8018 25616 -7958
rect 25676 -8018 25696 -7958
rect 25272 -8153 25372 -8152
rect 25267 -8251 25273 -8153
rect 25371 -8251 25377 -8153
rect 10604 -13353 10704 -13352
rect 10599 -13451 10605 -13353
rect 10703 -13451 10709 -13353
rect 10604 -13452 10704 -13451
rect 25272 -13586 25372 -8251
rect 25596 -13353 25696 -8018
rect 25591 -13451 25597 -13353
rect 25695 -13451 25701 -13353
rect 25596 -13452 25696 -13451
rect 25272 -13646 25300 -13586
rect 25360 -13646 25372 -13586
rect 25272 -13662 25372 -13646
rect 25402 -26153 25502 -26152
rect 40300 -26153 40400 -26152
rect 25397 -26251 25403 -26153
rect 25501 -26251 25507 -26153
rect 40295 -26251 40301 -26153
rect 40399 -26251 40405 -26153
rect 25402 -26252 25502 -26251
rect 40300 -26252 40400 -26251
<< via3 >>
rect 15532 3904 15914 4204
rect 23666 3904 24344 4204
rect 26114 3904 26714 4204
rect 30746 3904 31346 4204
rect 17600 3640 17696 3726
rect 18180 3640 18276 3726
rect 18780 3640 18876 3726
rect 19380 3640 19476 3726
rect 19980 3640 20076 3726
rect 20580 3640 20676 3726
rect 21180 3640 21276 3726
rect 21780 3640 21876 3726
rect 22380 3640 22476 3726
rect 26362 3640 26458 3726
rect 26942 3640 27038 3726
rect 27542 3640 27638 3726
rect 28142 3640 28238 3726
rect 28742 3640 28838 3726
rect 29342 3640 29438 3726
rect 29942 3640 30038 3726
rect 30542 3640 30638 3726
rect 31142 3640 31238 3726
rect 15532 -1552 15914 -1252
rect 23666 -1552 24344 -1252
rect 26114 -1552 26714 -1252
rect 30746 -1552 31346 -1252
rect 25273 -8251 25371 -8153
rect 10605 -13357 10703 -13353
rect 10605 -13447 10609 -13357
rect 10609 -13447 10699 -13357
rect 10699 -13447 10703 -13357
rect 10605 -13451 10703 -13447
rect 25597 -13451 25695 -13353
rect 25403 -26157 25501 -26153
rect 25403 -26247 25407 -26157
rect 25407 -26247 25497 -26157
rect 25497 -26247 25501 -26157
rect 25403 -26251 25501 -26247
rect 40301 -26157 40399 -26153
rect 40301 -26247 40305 -26157
rect 40305 -26247 40395 -26157
rect 40395 -26247 40399 -26157
rect 40301 -26251 40399 -26247
<< metal4 >>
rect 10584 4204 40288 4388
rect 10584 3904 15532 4204
rect 15914 3904 23666 4204
rect 24344 3904 26114 4204
rect 26714 3904 30746 4204
rect 31346 3904 40288 4204
rect 10584 3726 40288 3904
rect 10584 3640 17600 3726
rect 17696 3640 18180 3726
rect 18276 3640 18780 3726
rect 18876 3640 19380 3726
rect 19476 3640 19980 3726
rect 20076 3640 20580 3726
rect 20676 3640 21180 3726
rect 21276 3640 21780 3726
rect 21876 3640 22380 3726
rect 22476 3640 26362 3726
rect 26458 3640 26942 3726
rect 27038 3640 27542 3726
rect 27638 3640 28142 3726
rect 28238 3640 28742 3726
rect 28838 3640 29342 3726
rect 29438 3640 29942 3726
rect 30038 3640 30542 3726
rect 30638 3640 31142 3726
rect 31238 3640 40288 3726
rect 10584 3588 40288 3640
rect 15348 -940 31530 -936
rect 10744 -974 41209 -940
rect 10744 -1252 40432 -974
rect 10744 -1552 15532 -1252
rect 15914 -1552 23666 -1252
rect 24344 -1552 26114 -1252
rect 26714 -1552 30746 -1252
rect 31346 -1552 40432 -1252
rect 10744 -2722 40432 -1552
rect 41178 -2722 41209 -974
rect 10744 -2750 41209 -2722
rect 25158 -8153 25372 -8152
rect 25158 -8251 25273 -8153
rect 25371 -8251 25372 -8153
rect 25158 -8252 25372 -8251
rect 9780 -9856 12644 -9850
rect 24250 -9856 26734 -9850
rect 9780 -9878 40292 -9856
rect 9780 -11722 9814 -9878
rect 10548 -11722 40292 -9878
rect 9780 -11754 40292 -11722
rect 10604 -13353 10844 -13352
rect 10604 -13451 10605 -13353
rect 10703 -13451 10844 -13353
rect 10604 -13452 10844 -13451
rect 25596 -13353 25860 -13352
rect 25596 -13451 25597 -13353
rect 25695 -13451 25860 -13353
rect 25596 -13452 25860 -13451
rect 10740 -18880 41204 -18850
rect 10740 -20726 40432 -18880
rect 41166 -20726 41204 -18880
rect 10740 -20752 41204 -20726
rect 25190 -26153 25502 -26152
rect 25190 -26251 25403 -26153
rect 25501 -26251 25502 -26153
rect 25190 -26252 25502 -26251
rect 40190 -26153 40400 -26152
rect 40190 -26251 40301 -26153
rect 40399 -26251 40400 -26153
rect 40190 -26252 40400 -26251
rect 10586 -28650 11168 -27850
rect 24488 -28650 26804 -27850
<< via4 >>
rect 9784 3588 10584 4388
rect 40432 -2722 41178 -974
rect 9814 -11722 10548 -9878
rect 40432 -20726 41166 -18880
rect 9786 -28650 10586 -27850
<< metal5 >>
rect 9786 4412 10586 4472
rect 9760 4388 10608 4412
rect 9760 3588 9784 4388
rect 10584 3588 10608 4388
rect 9760 3564 10608 3588
rect 9786 -9878 10586 3564
rect 9786 -11722 9814 -9878
rect 10548 -11722 10586 -9878
rect 9786 -27826 10586 -11722
rect 40402 -974 41202 4472
rect 40402 -2722 40432 -974
rect 41178 -2722 41202 -974
rect 40402 -18880 41202 -2722
rect 40402 -20726 40432 -18880
rect 41166 -20726 41202 -18880
rect 9762 -27850 10610 -27826
rect 9762 -28650 9786 -27850
rect 10586 -28650 10610 -27850
rect 9762 -28674 10610 -28650
rect 9786 -28686 10586 -28674
rect 40402 -28686 41202 -20726
use cs_ring_osc_stage  cs_ring_osc_stage_2 cs_ring_osc_stage
timestamp 1623971255
transform 1 0 15840 0 1 -30350
box -5100 1696 9450 10400
use cs_ring_osc_stage  cs_ring_osc_stage_3
timestamp 1623971255
transform 1 0 30840 0 1 -30350
box -5100 1696 9450 10400
use cs_ring_osc_stage  cs_ring_osc_stage_1
timestamp 1623971255
transform -1 0 20194 0 -1 -9254
box -5100 1696 9450 10400
use cs_ring_osc_stage  cs_ring_osc_stage_4
timestamp 1623971255
transform -1 0 35194 0 -1 -9254
box -5100 1696 9450 10400
use cs_ring_osc_stage  cs_ring_osc_stage_0
timestamp 1623971255
transform 1 0 15840 0 1 -12350
box -5100 1696 9450 10400
use cs_ring_osc_stage  cs_ring_osc_stage_5
timestamp 1623971255
transform 1 0 30840 0 1 -12350
box -5100 1696 9450 10400
use sky130_fd_pr__nfet_01v8_V6PJ6N  sky130_fd_pr__nfet_01v8_V6PJ6N_0
timestamp 1623971255
transform 1 0 19941 0 -1 3144
box -2319 -188 2319 188
use sky130_fd_pr__pfet_01v8_hvt_GK2P2M  sky130_fd_pr__pfet_01v8_hvt_GK2P2M_0
timestamp 1623971255
transform 1 0 19941 0 -1 593
box -4187 -900 4187 900
use sky130_fd_pr__nfet_01v8_V6PJ6N  sky130_fd_pr__nfet_01v8_V6PJ6N_1
timestamp 1623971255
transform 1 0 28703 0 -1 3144
box -2319 -188 2319 188
use sky130_fd_pr__pfet_01v8_hvt_8Q5PU3  sky130_fd_pr__pfet_01v8_hvt_8Q5PU3_0
timestamp 1623971255
transform 1 0 28704 0 -1 1213
box -2355 -700 2355 700
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623971255
transform 1 0 31818 0 -1 2490
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623971255
transform 1 0 31542 0 -1 2490
box -38 -48 314 592
<< labels >>
flabel metal2 16596 1582 16604 1588 5 FreeSans 480 0 0 0 vpbias
flabel metal1 18498 3414 18504 3422 5 FreeSans 480 0 0 0 vctrl
flabel metal1 32398 2246 32414 2260 1 FreeSans 480 0 0 0 voscbuf
flabel metal1 31098 2304 31114 2316 1 FreeSans 480 0 0 0 vosc
flabel metal1 31796 2256 31804 2260 1 FreeSans 480 0 0 0 vosc2
flabel metal4 13612 3930 13632 3948 1 FreeSans 480 0 0 0 VSS
flabel metal4 13272 -1542 13284 -1524 1 FreeSans 480 0 0 0 VDD
<< properties >>
string FIXED_BBOX 20128 1902 25472 3682
<< end >>

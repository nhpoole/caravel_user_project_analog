magic
tech sky130A
magscale 1 2
timestamp 1624300568
<< nwell >>
rect -2454 122 3321 444
rect -2622 -634 3320 -398
rect -2622 -730 -2260 -634
rect -2242 -730 3320 -634
rect -2622 -966 3320 -730
rect -2622 -2054 3320 -1486
rect -2622 -2896 3320 -2574
<< pwell >>
rect -2582 -342 3280 66
rect -2582 -1430 3280 -1022
rect -2582 -2518 3280 -2110
<< locali >>
rect -2584 -155 -2555 -121
rect -2521 -155 -2492 -121
rect 3190 -155 3219 -121
rect 3253 -155 3282 -121
rect -2567 -198 -2509 -155
rect 3207 -198 3265 -155
rect -2567 -665 -2509 -622
rect 3207 -665 3265 -622
rect -2584 -699 -2555 -665
rect -2521 -699 -2492 -665
rect 3190 -699 3219 -665
rect 3253 -699 3282 -665
rect -2567 -742 -2509 -699
rect 3207 -742 3265 -699
rect -2567 -1209 -2509 -1166
rect 3207 -1209 3265 -1166
rect -2584 -1243 -2555 -1209
rect -2521 -1243 -2492 -1209
rect 3190 -1243 3219 -1209
rect 3253 -1243 3282 -1209
rect -2567 -1286 -2509 -1243
rect 3207 -1286 3265 -1243
rect -2567 -1753 -2509 -1710
rect 3207 -1753 3265 -1710
rect -2584 -1787 -2555 -1753
rect -2521 -1787 -2492 -1753
rect 3190 -1787 3219 -1753
rect 3253 -1787 3282 -1753
rect -2567 -1830 -2509 -1787
rect 3207 -1830 3265 -1787
rect -2567 -2297 -2509 -2254
rect 3207 -2297 3265 -2254
rect -2584 -2331 -2555 -2297
rect -2521 -2331 -2492 -2297
rect 3190 -2331 3219 -2297
rect 3253 -2331 3282 -2297
rect -2567 -2374 -2509 -2331
rect 3207 -2374 3265 -2331
rect -2567 -2841 -2509 -2798
rect 3207 -2841 3265 -2798
rect -2584 -2875 -2555 -2841
rect -2521 -2875 -2492 -2841
rect 3190 -2875 3219 -2841
rect 3253 -2875 3282 -2841
<< viali >>
rect -2214 98 -2166 146
rect -1962 40 -1914 88
rect -552 78 -504 126
rect -436 78 -388 126
rect -324 78 -276 126
rect -192 78 -144 126
rect -82 78 -34 126
rect 34 78 82 126
rect 166 76 214 124
rect -858 -40 -810 8
rect -2555 -155 -2521 -121
rect 3219 -155 3253 -121
rect 1842 -288 1890 -240
rect -1962 -364 -1914 -316
rect -2218 -412 -2170 -364
rect -552 -402 -504 -354
rect -436 -402 -388 -354
rect -324 -402 -276 -354
rect -192 -402 -144 -354
rect -82 -402 -34 -354
rect 34 -402 82 -354
rect 170 -400 218 -352
rect 736 -364 784 -316
rect 2146 -402 2194 -354
rect 2262 -402 2310 -354
rect 2374 -402 2422 -354
rect 2506 -402 2554 -354
rect 2616 -402 2664 -354
rect 2732 -402 2780 -354
rect 2864 -400 2912 -352
rect 480 -454 528 -406
rect -858 -586 -810 -538
rect -2555 -699 -2521 -665
rect 3219 -699 3253 -665
rect 1840 -826 1888 -778
rect -2218 -958 -2170 -910
rect -1962 -1048 -1914 -1000
rect -552 -1010 -504 -962
rect -436 -1010 -388 -962
rect -324 -1010 -276 -962
rect -192 -1010 -144 -962
rect -82 -1010 -34 -962
rect 34 -1010 82 -962
rect 166 -1012 218 -964
rect 480 -998 528 -950
rect 736 -1048 784 -1000
rect 2146 -1010 2194 -962
rect 2262 -1010 2310 -962
rect 2374 -1010 2422 -962
rect 2506 -1010 2554 -962
rect 2616 -1010 2664 -962
rect 2732 -1010 2780 -962
rect 2864 -1012 2912 -964
rect -858 -1130 -810 -1082
rect -2555 -1243 -2521 -1209
rect 3219 -1243 3253 -1209
rect 1840 -1370 1888 -1322
rect -1962 -1452 -1914 -1404
rect -2218 -1502 -2170 -1454
rect -552 -1490 -504 -1442
rect -436 -1490 -388 -1442
rect -324 -1490 -276 -1442
rect -192 -1490 -144 -1442
rect -82 -1490 -34 -1442
rect 34 -1490 82 -1442
rect 166 -1488 214 -1440
rect 736 -1452 784 -1404
rect 2146 -1490 2194 -1442
rect 2262 -1490 2310 -1442
rect 2374 -1490 2422 -1442
rect 2506 -1490 2554 -1442
rect 2616 -1490 2664 -1442
rect 2732 -1490 2780 -1442
rect 2864 -1488 2916 -1440
rect 480 -1542 528 -1494
rect -858 -1674 -810 -1626
rect -2555 -1787 -2521 -1753
rect 3219 -1787 3253 -1753
rect 1840 -1914 1888 -1866
rect -2218 -2046 -2170 -1998
rect -1962 -2136 -1914 -2088
rect -552 -2098 -504 -2050
rect -436 -2098 -388 -2050
rect -324 -2098 -276 -2050
rect -192 -2098 -144 -2050
rect -82 -2098 -34 -2050
rect 34 -2098 82 -2050
rect 166 -2100 214 -2052
rect 480 -2088 528 -2040
rect 736 -2136 784 -2088
rect 2146 -2098 2194 -2050
rect 2262 -2098 2310 -2050
rect 2374 -2098 2422 -2050
rect 2506 -2098 2554 -2050
rect 2616 -2098 2664 -2050
rect 2732 -2098 2780 -2050
rect 2868 -2100 2916 -2052
rect -858 -2216 -810 -2168
rect -2555 -2331 -2521 -2297
rect 3219 -2331 3253 -2297
rect 1840 -2460 1888 -2412
rect -1962 -2540 -1914 -2492
rect -2218 -2588 -2170 -2540
rect -552 -2578 -504 -2530
rect -436 -2578 -388 -2530
rect -324 -2578 -276 -2530
rect -192 -2578 -144 -2530
rect -82 -2578 -34 -2530
rect 34 -2578 82 -2530
rect 166 -2576 218 -2528
rect 488 -2570 536 -2522
rect 736 -2540 784 -2492
rect 2146 -2578 2194 -2530
rect 2262 -2578 2310 -2530
rect 2374 -2578 2422 -2530
rect 2506 -2578 2554 -2530
rect 2616 -2578 2664 -2530
rect 2732 -2578 2780 -2530
rect 2864 -2576 2912 -2528
rect -858 -2760 -810 -2712
rect -2555 -2875 -2521 -2841
rect 3219 -2875 3253 -2841
<< metal1 >>
rect -2492 358 -2242 454
rect 242 442 3190 454
rect 242 370 292 442
rect 388 370 3190 442
rect 242 358 3190 370
rect -2674 146 -2154 152
rect -2674 98 -2214 146
rect -2166 98 -2154 146
rect -564 126 -376 132
rect -2674 92 -2154 98
rect -1968 94 -1908 100
rect -1974 34 -1968 94
rect -1908 34 -1902 94
rect -564 78 -552 126
rect -504 78 -436 126
rect -388 78 -376 126
rect -564 72 -376 78
rect -336 126 94 132
rect 160 130 220 136
rect -336 78 -324 126
rect -276 78 -192 126
rect -144 78 -82 126
rect -34 78 34 126
rect 82 78 94 126
rect -336 72 94 78
rect 154 70 160 130
rect 220 70 226 130
rect 160 64 220 70
rect -1968 28 -1908 34
rect -864 14 -804 20
rect -870 -46 -864 14
rect -804 -46 -798 14
rect -864 -52 -804 -46
rect -2584 -102 -2242 -90
rect -2584 -121 -2388 -102
rect -2584 -155 -2555 -121
rect -2521 -155 -2388 -121
rect -2584 -174 -2388 -155
rect -2292 -174 -2242 -102
rect -2584 -186 -2242 -174
rect 242 -186 456 -90
rect 2938 -102 3282 -90
rect 2938 -174 2990 -102
rect 3086 -121 3282 -102
rect 3086 -155 3219 -121
rect 3253 -155 3282 -121
rect 3086 -174 3282 -155
rect 2938 -186 3282 -174
rect 1836 -234 1896 -228
rect 1830 -294 1836 -234
rect 1896 -294 1902 -234
rect 1836 -300 1896 -294
rect -1968 -310 -1908 -304
rect 730 -310 790 -304
rect -2224 -358 -2164 -352
rect -2230 -418 -2224 -358
rect -2164 -418 -2158 -358
rect -1974 -370 -1968 -310
rect -1908 -370 -1902 -310
rect -564 -354 -376 -348
rect -1968 -376 -1908 -370
rect -564 -402 -552 -354
rect -504 -402 -436 -354
rect -388 -402 -376 -354
rect -564 -408 -376 -402
rect -336 -354 94 -348
rect -336 -402 -324 -354
rect -276 -402 -192 -354
rect -144 -402 -82 -354
rect -34 -402 34 -354
rect 82 -402 94 -354
rect -336 -408 94 -402
rect 152 -406 158 -346
rect 218 -406 230 -346
rect 724 -370 730 -310
rect 790 -370 796 -310
rect 2858 -346 2918 -340
rect 2134 -354 2322 -348
rect 730 -376 790 -370
rect 474 -400 534 -394
rect -2224 -424 -2164 -418
rect 468 -460 474 -400
rect 534 -460 540 -400
rect 2134 -402 2146 -354
rect 2194 -402 2262 -354
rect 2310 -402 2322 -354
rect 2134 -408 2322 -402
rect 2362 -354 2792 -348
rect 2362 -402 2374 -354
rect 2422 -402 2506 -354
rect 2554 -402 2616 -354
rect 2664 -402 2732 -354
rect 2780 -402 2792 -354
rect 2362 -408 2792 -402
rect 2852 -406 2858 -346
rect 2918 -406 2924 -346
rect 2858 -412 2918 -406
rect 474 -466 534 -460
rect -864 -532 -804 -526
rect -870 -592 -864 -532
rect -804 -592 -798 -532
rect -864 -598 -804 -592
rect -2584 -665 -2242 -634
rect -2584 -699 -2555 -665
rect -2521 -699 -2242 -665
rect -2584 -730 -2242 -699
rect 242 -646 456 -634
rect 242 -718 292 -646
rect 388 -718 456 -646
rect 242 -730 456 -718
rect 2936 -665 3282 -634
rect 2936 -699 3219 -665
rect 3253 -699 3282 -665
rect 2936 -730 3282 -699
rect 1834 -772 1894 -766
rect 1828 -832 1834 -772
rect 1894 -832 1900 -772
rect 1834 -838 1894 -832
rect -2224 -904 -2164 -898
rect -2230 -964 -2224 -904
rect -2164 -964 -2158 -904
rect 474 -944 534 -938
rect -564 -962 -376 -956
rect -2224 -970 -2164 -964
rect -1968 -994 -1908 -988
rect -1974 -1054 -1968 -994
rect -1908 -1054 -1902 -994
rect -564 -1010 -552 -962
rect -504 -1010 -436 -962
rect -388 -1010 -376 -962
rect -564 -1016 -376 -1010
rect -336 -962 94 -956
rect 160 -958 220 -952
rect -336 -1010 -324 -962
rect -276 -1010 -192 -962
rect -144 -1010 -82 -962
rect -34 -1010 34 -962
rect 82 -1010 94 -962
rect -336 -1016 94 -1010
rect 154 -1018 160 -958
rect 220 -1018 226 -958
rect 468 -1004 474 -944
rect 534 -1004 540 -944
rect 2134 -962 2322 -956
rect 730 -994 790 -988
rect 474 -1010 534 -1004
rect 160 -1024 220 -1018
rect 724 -1054 730 -994
rect 790 -1054 796 -994
rect 2134 -1010 2146 -962
rect 2194 -1010 2262 -962
rect 2310 -1010 2322 -962
rect 2134 -1016 2322 -1010
rect 2362 -962 2792 -956
rect 2858 -958 2918 -952
rect 2362 -1010 2374 -962
rect 2422 -1010 2506 -962
rect 2554 -1010 2616 -962
rect 2664 -1010 2732 -962
rect 2780 -1010 2792 -962
rect 2362 -1016 2792 -1010
rect 2852 -1018 2858 -958
rect 2918 -1018 2924 -958
rect 2858 -1024 2918 -1018
rect -1968 -1060 -1908 -1054
rect 730 -1060 790 -1054
rect -864 -1076 -804 -1070
rect -870 -1136 -864 -1076
rect -804 -1136 -798 -1076
rect -864 -1142 -804 -1136
rect -2584 -1190 -2224 -1178
rect -2584 -1209 -2388 -1190
rect -2584 -1243 -2555 -1209
rect -2521 -1243 -2388 -1209
rect -2584 -1262 -2388 -1243
rect -2292 -1262 -2224 -1190
rect -2584 -1274 -2224 -1262
rect 242 -1274 456 -1178
rect 2938 -1190 3282 -1178
rect 2938 -1262 2990 -1190
rect 3086 -1209 3282 -1190
rect 3086 -1243 3219 -1209
rect 3253 -1243 3282 -1209
rect 3086 -1262 3282 -1243
rect 2938 -1274 3282 -1262
rect 1834 -1316 1894 -1310
rect 1828 -1376 1834 -1316
rect 1894 -1376 1900 -1316
rect 1834 -1382 1894 -1376
rect -1968 -1398 -1908 -1392
rect 730 -1398 790 -1392
rect -2224 -1448 -2164 -1442
rect -2230 -1508 -2224 -1448
rect -2164 -1508 -2158 -1448
rect -1974 -1458 -1968 -1398
rect -1908 -1458 -1902 -1398
rect 160 -1434 220 -1428
rect -564 -1442 -376 -1436
rect -1968 -1464 -1908 -1458
rect -564 -1490 -552 -1442
rect -504 -1490 -436 -1442
rect -388 -1490 -376 -1442
rect -564 -1496 -376 -1490
rect -336 -1442 94 -1436
rect -336 -1490 -324 -1442
rect -276 -1490 -192 -1442
rect -144 -1490 -82 -1442
rect -34 -1490 34 -1442
rect 82 -1490 94 -1442
rect -336 -1496 94 -1490
rect 154 -1494 160 -1434
rect 220 -1494 226 -1434
rect 724 -1458 730 -1398
rect 790 -1458 796 -1398
rect 2858 -1434 2918 -1428
rect 2134 -1442 2322 -1436
rect 730 -1464 790 -1458
rect 474 -1488 534 -1482
rect 160 -1500 220 -1494
rect -2224 -1514 -2164 -1508
rect 468 -1548 474 -1488
rect 534 -1548 540 -1488
rect 2134 -1490 2146 -1442
rect 2194 -1490 2262 -1442
rect 2310 -1490 2322 -1442
rect 2134 -1496 2322 -1490
rect 2362 -1442 2792 -1436
rect 2362 -1490 2374 -1442
rect 2422 -1490 2506 -1442
rect 2554 -1490 2616 -1442
rect 2664 -1490 2732 -1442
rect 2780 -1490 2792 -1442
rect 2362 -1496 2792 -1490
rect 2852 -1494 2858 -1434
rect 2918 -1494 2924 -1434
rect 2858 -1500 2918 -1494
rect 474 -1554 534 -1548
rect -864 -1620 -804 -1614
rect -870 -1680 -864 -1620
rect -804 -1680 -798 -1620
rect -864 -1686 -804 -1680
rect -2584 -1753 -2242 -1722
rect -2584 -1787 -2555 -1753
rect -2521 -1787 -2242 -1753
rect -2584 -1818 -2242 -1787
rect 242 -1734 456 -1722
rect 242 -1806 292 -1734
rect 388 -1806 456 -1734
rect 242 -1818 456 -1806
rect 2936 -1753 3282 -1722
rect 2936 -1787 3219 -1753
rect 3253 -1787 3282 -1753
rect 2936 -1818 3282 -1787
rect 1834 -1860 1894 -1854
rect 1828 -1920 1834 -1860
rect 1894 -1920 1900 -1860
rect 1834 -1926 1894 -1920
rect -2224 -1992 -2164 -1986
rect -2230 -2052 -2224 -1992
rect -2164 -2052 -2158 -1992
rect 474 -2034 534 -2028
rect -564 -2050 -376 -2044
rect -2224 -2058 -2164 -2052
rect -1968 -2082 -1908 -2076
rect -1974 -2142 -1968 -2082
rect -1908 -2142 -1902 -2082
rect -564 -2098 -552 -2050
rect -504 -2098 -436 -2050
rect -388 -2098 -376 -2050
rect -564 -2104 -376 -2098
rect -336 -2050 94 -2044
rect 160 -2046 220 -2040
rect -336 -2098 -324 -2050
rect -276 -2098 -192 -2050
rect -144 -2098 -82 -2050
rect -34 -2098 34 -2050
rect 82 -2098 94 -2050
rect -336 -2104 94 -2098
rect 154 -2106 160 -2046
rect 220 -2106 226 -2046
rect 468 -2094 474 -2034
rect 534 -2094 540 -2034
rect 2134 -2050 2322 -2044
rect 730 -2082 790 -2076
rect 474 -2100 534 -2094
rect 160 -2112 220 -2106
rect 724 -2142 730 -2082
rect 790 -2142 796 -2082
rect 2134 -2098 2146 -2050
rect 2194 -2098 2262 -2050
rect 2310 -2098 2322 -2050
rect 2134 -2104 2322 -2098
rect 2362 -2050 2792 -2044
rect 2362 -2098 2374 -2050
rect 2422 -2098 2506 -2050
rect 2554 -2098 2616 -2050
rect 2664 -2098 2732 -2050
rect 2780 -2098 2792 -2050
rect 2362 -2104 2792 -2098
rect 2850 -2106 2856 -2046
rect 2916 -2106 2928 -2046
rect -1968 -2148 -1908 -2142
rect 730 -2148 790 -2142
rect -864 -2162 -804 -2156
rect -870 -2222 -864 -2162
rect -804 -2222 -798 -2162
rect -864 -2228 -804 -2222
rect -2584 -2278 -2224 -2266
rect -2584 -2297 -2388 -2278
rect -2584 -2331 -2555 -2297
rect -2521 -2331 -2388 -2297
rect -2584 -2350 -2388 -2331
rect -2292 -2350 -2224 -2278
rect -2584 -2362 -2224 -2350
rect 242 -2362 456 -2266
rect 2936 -2278 3282 -2266
rect 2936 -2350 2990 -2278
rect 3086 -2297 3282 -2278
rect 3086 -2331 3219 -2297
rect 3253 -2331 3282 -2297
rect 3086 -2350 3282 -2331
rect 2936 -2362 3282 -2350
rect 1834 -2406 1894 -2400
rect 1828 -2466 1834 -2406
rect 1894 -2466 1900 -2406
rect 1834 -2472 1894 -2466
rect -1968 -2486 -1908 -2480
rect 730 -2486 790 -2480
rect -2224 -2534 -2164 -2528
rect -2230 -2594 -2224 -2534
rect -2164 -2594 -2158 -2534
rect -1974 -2546 -1968 -2486
rect -1908 -2546 -1902 -2486
rect 482 -2516 542 -2510
rect 160 -2522 220 -2516
rect -564 -2530 -376 -2524
rect -1968 -2552 -1908 -2546
rect -564 -2578 -552 -2530
rect -504 -2578 -436 -2530
rect -388 -2578 -376 -2530
rect -564 -2584 -376 -2578
rect -336 -2530 94 -2524
rect -336 -2578 -324 -2530
rect -276 -2578 -192 -2530
rect -144 -2578 -82 -2530
rect -34 -2578 34 -2530
rect 82 -2578 94 -2530
rect -336 -2584 94 -2578
rect 154 -2582 160 -2522
rect 220 -2582 226 -2522
rect 476 -2576 482 -2516
rect 542 -2576 548 -2516
rect 724 -2546 730 -2486
rect 790 -2546 796 -2486
rect 2858 -2522 2918 -2516
rect 2134 -2530 2322 -2524
rect 730 -2552 790 -2546
rect 482 -2582 542 -2576
rect 2134 -2578 2146 -2530
rect 2194 -2578 2262 -2530
rect 2310 -2578 2322 -2530
rect 160 -2588 220 -2582
rect 2134 -2584 2322 -2578
rect 2362 -2530 2792 -2524
rect 2362 -2578 2374 -2530
rect 2422 -2578 2506 -2530
rect 2554 -2578 2616 -2530
rect 2664 -2578 2732 -2530
rect 2780 -2578 2792 -2530
rect 2362 -2584 2792 -2578
rect 2852 -2582 2858 -2522
rect 2918 -2582 2924 -2522
rect 2858 -2588 2918 -2582
rect -2224 -2600 -2164 -2594
rect -864 -2706 -804 -2700
rect -870 -2766 -864 -2706
rect -804 -2766 -798 -2706
rect -864 -2772 -804 -2766
rect -2584 -2841 -2242 -2810
rect -2584 -2875 -2555 -2841
rect -2521 -2875 -2242 -2841
rect -2584 -2906 -2242 -2875
rect 242 -2822 456 -2810
rect 242 -2894 292 -2822
rect 388 -2894 456 -2822
rect 242 -2906 456 -2894
rect 2936 -2841 3282 -2810
rect 2936 -2875 3219 -2841
rect 3253 -2875 3282 -2841
rect 2936 -2906 3282 -2875
<< via1 >>
rect 292 370 388 442
rect -1968 88 -1908 94
rect -1968 40 -1962 88
rect -1962 40 -1914 88
rect -1914 40 -1908 88
rect -1968 34 -1908 40
rect 160 124 220 130
rect 160 76 166 124
rect 166 76 214 124
rect 214 76 220 124
rect 160 70 220 76
rect -864 8 -804 14
rect -864 -40 -858 8
rect -858 -40 -810 8
rect -810 -40 -804 8
rect -864 -46 -804 -40
rect -2388 -174 -2292 -102
rect 2990 -174 3086 -102
rect 1836 -240 1896 -234
rect 1836 -288 1842 -240
rect 1842 -288 1890 -240
rect 1890 -288 1896 -240
rect 1836 -294 1896 -288
rect -2224 -364 -2164 -358
rect -2224 -412 -2218 -364
rect -2218 -412 -2170 -364
rect -2170 -412 -2164 -364
rect -2224 -418 -2164 -412
rect -1968 -316 -1908 -310
rect -1968 -364 -1962 -316
rect -1962 -364 -1914 -316
rect -1914 -364 -1908 -316
rect -1968 -370 -1908 -364
rect 158 -352 218 -346
rect 158 -400 170 -352
rect 170 -400 218 -352
rect 158 -406 218 -400
rect 730 -316 790 -310
rect 730 -364 736 -316
rect 736 -364 784 -316
rect 784 -364 790 -316
rect 730 -370 790 -364
rect 474 -406 534 -400
rect 474 -454 480 -406
rect 480 -454 528 -406
rect 528 -454 534 -406
rect 474 -460 534 -454
rect 2858 -352 2918 -346
rect 2858 -400 2864 -352
rect 2864 -400 2912 -352
rect 2912 -400 2918 -352
rect 2858 -406 2918 -400
rect -864 -538 -804 -532
rect -864 -586 -858 -538
rect -858 -586 -810 -538
rect -810 -586 -804 -538
rect -864 -592 -804 -586
rect 292 -718 388 -646
rect 1834 -778 1894 -772
rect 1834 -826 1840 -778
rect 1840 -826 1888 -778
rect 1888 -826 1894 -778
rect 1834 -832 1894 -826
rect -2224 -910 -2164 -904
rect -2224 -958 -2218 -910
rect -2218 -958 -2170 -910
rect -2170 -958 -2164 -910
rect -2224 -964 -2164 -958
rect -1968 -1000 -1908 -994
rect -1968 -1048 -1962 -1000
rect -1962 -1048 -1914 -1000
rect -1914 -1048 -1908 -1000
rect -1968 -1054 -1908 -1048
rect 160 -964 220 -958
rect 160 -1012 166 -964
rect 166 -1012 218 -964
rect 218 -1012 220 -964
rect 160 -1018 220 -1012
rect 474 -950 534 -944
rect 474 -998 480 -950
rect 480 -998 528 -950
rect 528 -998 534 -950
rect 474 -1004 534 -998
rect 730 -1000 790 -994
rect 730 -1048 736 -1000
rect 736 -1048 784 -1000
rect 784 -1048 790 -1000
rect 730 -1054 790 -1048
rect 2858 -964 2918 -958
rect 2858 -1012 2864 -964
rect 2864 -1012 2912 -964
rect 2912 -1012 2918 -964
rect 2858 -1018 2918 -1012
rect -864 -1082 -804 -1076
rect -864 -1130 -858 -1082
rect -858 -1130 -810 -1082
rect -810 -1130 -804 -1082
rect -864 -1136 -804 -1130
rect -2388 -1262 -2292 -1190
rect 2990 -1262 3086 -1190
rect 1834 -1322 1894 -1316
rect 1834 -1370 1840 -1322
rect 1840 -1370 1888 -1322
rect 1888 -1370 1894 -1322
rect 1834 -1376 1894 -1370
rect -2224 -1454 -2164 -1448
rect -2224 -1502 -2218 -1454
rect -2218 -1502 -2170 -1454
rect -2170 -1502 -2164 -1454
rect -2224 -1508 -2164 -1502
rect -1968 -1404 -1908 -1398
rect -1968 -1452 -1962 -1404
rect -1962 -1452 -1914 -1404
rect -1914 -1452 -1908 -1404
rect -1968 -1458 -1908 -1452
rect 160 -1440 220 -1434
rect 160 -1488 166 -1440
rect 166 -1488 214 -1440
rect 214 -1488 220 -1440
rect 160 -1494 220 -1488
rect 730 -1404 790 -1398
rect 730 -1452 736 -1404
rect 736 -1452 784 -1404
rect 784 -1452 790 -1404
rect 730 -1458 790 -1452
rect 474 -1494 534 -1488
rect 474 -1542 480 -1494
rect 480 -1542 528 -1494
rect 528 -1542 534 -1494
rect 474 -1548 534 -1542
rect 2858 -1440 2918 -1434
rect 2858 -1488 2864 -1440
rect 2864 -1488 2916 -1440
rect 2916 -1488 2918 -1440
rect 2858 -1494 2918 -1488
rect -864 -1626 -804 -1620
rect -864 -1674 -858 -1626
rect -858 -1674 -810 -1626
rect -810 -1674 -804 -1626
rect -864 -1680 -804 -1674
rect 292 -1806 388 -1734
rect 1834 -1866 1894 -1860
rect 1834 -1914 1840 -1866
rect 1840 -1914 1888 -1866
rect 1888 -1914 1894 -1866
rect 1834 -1920 1894 -1914
rect -2224 -1998 -2164 -1992
rect -2224 -2046 -2218 -1998
rect -2218 -2046 -2170 -1998
rect -2170 -2046 -2164 -1998
rect -2224 -2052 -2164 -2046
rect -1968 -2088 -1908 -2082
rect -1968 -2136 -1962 -2088
rect -1962 -2136 -1914 -2088
rect -1914 -2136 -1908 -2088
rect -1968 -2142 -1908 -2136
rect 160 -2052 220 -2046
rect 160 -2100 166 -2052
rect 166 -2100 214 -2052
rect 214 -2100 220 -2052
rect 160 -2106 220 -2100
rect 474 -2040 534 -2034
rect 474 -2088 480 -2040
rect 480 -2088 528 -2040
rect 528 -2088 534 -2040
rect 474 -2094 534 -2088
rect 730 -2088 790 -2082
rect 730 -2136 736 -2088
rect 736 -2136 784 -2088
rect 784 -2136 790 -2088
rect 730 -2142 790 -2136
rect 2856 -2052 2916 -2046
rect 2856 -2100 2868 -2052
rect 2868 -2100 2916 -2052
rect 2856 -2106 2916 -2100
rect -864 -2168 -804 -2162
rect -864 -2216 -858 -2168
rect -858 -2216 -810 -2168
rect -810 -2216 -804 -2168
rect -864 -2222 -804 -2216
rect -2388 -2350 -2292 -2278
rect 2990 -2350 3086 -2278
rect 1834 -2412 1894 -2406
rect 1834 -2460 1840 -2412
rect 1840 -2460 1888 -2412
rect 1888 -2460 1894 -2412
rect 1834 -2466 1894 -2460
rect -2224 -2540 -2164 -2534
rect -2224 -2588 -2218 -2540
rect -2218 -2588 -2170 -2540
rect -2170 -2588 -2164 -2540
rect -2224 -2594 -2164 -2588
rect -1968 -2492 -1908 -2486
rect -1968 -2540 -1962 -2492
rect -1962 -2540 -1914 -2492
rect -1914 -2540 -1908 -2492
rect -1968 -2546 -1908 -2540
rect 160 -2528 220 -2522
rect 160 -2576 166 -2528
rect 166 -2576 218 -2528
rect 218 -2576 220 -2528
rect 160 -2582 220 -2576
rect 482 -2522 542 -2516
rect 482 -2570 488 -2522
rect 488 -2570 536 -2522
rect 536 -2570 542 -2522
rect 482 -2576 542 -2570
rect 730 -2492 790 -2486
rect 730 -2540 736 -2492
rect 736 -2540 784 -2492
rect 784 -2540 790 -2492
rect 730 -2546 790 -2540
rect 2858 -2528 2918 -2522
rect 2858 -2576 2864 -2528
rect 2864 -2576 2912 -2528
rect 2912 -2576 2918 -2528
rect 2858 -2582 2918 -2576
rect -864 -2712 -804 -2706
rect -864 -2760 -858 -2712
rect -858 -2760 -810 -2712
rect -810 -2760 -804 -2712
rect -864 -2766 -804 -2760
rect 292 -2894 388 -2822
<< metal2 >>
rect 280 442 400 454
rect 280 370 292 442
rect 388 370 400 442
rect 280 358 400 370
rect -1968 94 160 130
rect -1908 70 160 94
rect 220 70 226 130
rect -1968 28 -1908 34
rect -864 14 -804 20
rect -2400 -102 -2280 -90
rect -2400 -174 -2388 -102
rect -2292 -174 -2280 -102
rect -864 -106 -804 -46
rect -2400 -186 -2280 -174
rect -2224 -166 -804 -106
rect -2224 -358 -2164 -166
rect 1836 -234 1896 104
rect 2978 -102 3098 -90
rect 2978 -174 2990 -102
rect 3086 -174 3098 -102
rect 2978 -186 3098 -174
rect 1830 -294 1836 -234
rect 1896 -294 1902 -234
rect -1968 -310 -1908 -304
rect 730 -310 790 -304
rect 158 -346 224 -340
rect -1908 -370 158 -346
rect -1968 -406 158 -370
rect 218 -406 224 -346
rect 790 -370 2858 -346
rect 158 -412 224 -406
rect 474 -400 534 -394
rect -2224 -424 -2164 -418
rect 730 -406 2858 -370
rect 2918 -406 2924 -346
rect -864 -532 -804 -526
rect -864 -652 -804 -592
rect -2224 -712 -804 -652
rect 280 -646 400 -634
rect -2224 -904 -2164 -712
rect 280 -718 292 -646
rect 388 -718 400 -646
rect 474 -652 534 -460
rect 474 -712 1894 -652
rect 280 -730 400 -718
rect 1834 -772 1894 -712
rect 1834 -838 1894 -832
rect 474 -944 534 -938
rect -2224 -970 -2164 -964
rect -1968 -994 160 -958
rect -1908 -1018 160 -994
rect 220 -1018 226 -958
rect -1968 -1060 -1908 -1054
rect -864 -1076 -804 -1070
rect -2400 -1190 -2280 -1178
rect -2400 -1262 -2388 -1190
rect -2292 -1262 -2280 -1190
rect -864 -1196 -804 -1136
rect -2400 -1274 -2280 -1262
rect -2224 -1256 -804 -1196
rect 474 -1196 534 -1004
rect 730 -994 2858 -958
rect 790 -1018 2858 -994
rect 2918 -1018 2924 -958
rect 730 -1060 790 -1054
rect 2978 -1190 3098 -1178
rect 474 -1256 1894 -1196
rect -2224 -1448 -2164 -1256
rect 1834 -1316 1894 -1256
rect 2978 -1262 2990 -1190
rect 3086 -1262 3098 -1190
rect 2978 -1274 3098 -1262
rect 1834 -1382 1894 -1376
rect -1968 -1398 -1908 -1392
rect 730 -1398 790 -1392
rect -1908 -1458 160 -1434
rect -1968 -1494 160 -1458
rect 220 -1494 226 -1434
rect 790 -1458 2858 -1434
rect 474 -1488 534 -1482
rect -2224 -1514 -2164 -1508
rect 730 -1494 2858 -1458
rect 2918 -1494 2924 -1434
rect -864 -1620 -804 -1614
rect -864 -1740 -804 -1680
rect -2224 -1800 -804 -1740
rect 280 -1734 400 -1722
rect -2224 -1992 -2164 -1800
rect 280 -1806 292 -1734
rect 388 -1806 400 -1734
rect 474 -1740 534 -1548
rect 474 -1800 1894 -1740
rect 280 -1818 400 -1806
rect 1834 -1860 1894 -1800
rect 1834 -1926 1894 -1920
rect 474 -2034 534 -2028
rect -2224 -2058 -2164 -2052
rect -1968 -2082 160 -2046
rect -1908 -2106 160 -2082
rect 220 -2106 226 -2046
rect 2856 -2046 2922 -2040
rect -1968 -2148 -1908 -2142
rect -864 -2162 -804 -2156
rect -2400 -2278 -2280 -2266
rect -2400 -2350 -2388 -2278
rect -2292 -2350 -2280 -2278
rect -864 -2282 -804 -2222
rect -2400 -2362 -2280 -2350
rect -2224 -2342 -804 -2282
rect 474 -2286 534 -2094
rect 730 -2082 2856 -2046
rect 790 -2106 2856 -2082
rect 2916 -2106 2922 -2046
rect 2856 -2112 2922 -2106
rect 730 -2148 790 -2142
rect 2978 -2278 3098 -2266
rect -2224 -2534 -2164 -2342
rect 474 -2346 1894 -2286
rect 1834 -2406 1894 -2346
rect 2978 -2350 2990 -2278
rect 3086 -2350 3098 -2278
rect 2978 -2362 3098 -2350
rect 1834 -2472 1894 -2466
rect -1968 -2486 -1908 -2480
rect 730 -2486 790 -2480
rect 482 -2516 542 -2510
rect -1908 -2546 160 -2522
rect -1968 -2582 160 -2546
rect 220 -2582 226 -2522
rect 376 -2576 482 -2516
rect -2224 -2600 -2164 -2594
rect -864 -2706 -804 -2700
rect 376 -2706 436 -2576
rect 482 -2582 542 -2576
rect 790 -2546 2858 -2522
rect 730 -2582 2858 -2546
rect 2918 -2582 2924 -2522
rect -804 -2766 436 -2706
rect -864 -2772 -804 -2766
rect 280 -2822 400 -2810
rect 280 -2894 292 -2822
rect 388 -2894 400 -2822
rect 280 -2906 400 -2894
<< via2 >>
rect 292 370 388 442
rect -2388 -174 -2292 -102
rect 2990 -174 3086 -102
rect 292 -718 388 -646
rect -2388 -1262 -2292 -1190
rect 2990 -1262 3086 -1190
rect 292 -1806 388 -1734
rect -2388 -2350 -2292 -2278
rect 2990 -2350 3086 -2278
rect 292 -2894 388 -2822
<< metal3 >>
rect 280 442 400 454
rect 280 370 292 442
rect 388 370 400 442
rect 280 358 400 370
rect -2400 -102 -2280 -90
rect -2400 -174 -2388 -102
rect -2292 -174 -2280 -102
rect -2400 -186 -2280 -174
rect 2978 -102 3098 -90
rect 2978 -174 2990 -102
rect 3086 -174 3098 -102
rect 2978 -186 3098 -174
rect 280 -646 400 -634
rect 280 -718 292 -646
rect 388 -718 400 -646
rect 280 -730 400 -718
rect -2400 -1190 -2280 -1178
rect -2400 -1262 -2388 -1190
rect -2292 -1262 -2280 -1190
rect -2400 -1274 -2280 -1262
rect 2978 -1190 3098 -1178
rect 2978 -1262 2990 -1190
rect 3086 -1262 3098 -1190
rect 2978 -1274 3098 -1262
rect 280 -1734 400 -1722
rect 280 -1806 292 -1734
rect 388 -1806 400 -1734
rect 280 -1818 400 -1806
rect -2400 -2278 -2280 -2266
rect -2400 -2350 -2388 -2278
rect -2292 -2350 -2280 -2278
rect -2400 -2362 -2280 -2350
rect 2978 -2278 3098 -2266
rect 2978 -2350 2990 -2278
rect 3086 -2350 3098 -2278
rect 2978 -2362 3098 -2350
rect 280 -2822 400 -2810
rect 280 -2894 292 -2822
rect 388 -2894 400 -2822
rect 280 -2906 400 -2894
<< via3 >>
rect 292 370 388 442
rect -2388 -174 -2292 -102
rect 2990 -174 3086 -102
rect 292 -718 388 -646
rect -2388 -1262 -2292 -1190
rect 2990 -1262 3086 -1190
rect 292 -1806 388 -1734
rect -2388 -2350 -2292 -2278
rect 2990 -2350 3086 -2278
rect 292 -2894 388 -2822
<< metal4 >>
rect -2400 -102 -2280 454
rect -2400 -174 -2388 -102
rect -2292 -174 -2280 -102
rect -2400 -1190 -2280 -174
rect -2400 -1262 -2388 -1190
rect -2292 -1262 -2280 -1190
rect -2400 -2278 -2280 -1262
rect -2400 -2350 -2388 -2278
rect -2292 -2350 -2280 -2278
rect -2400 -2906 -2280 -2350
rect 280 442 400 454
rect 280 370 292 442
rect 388 370 400 442
rect 280 -646 400 370
rect 280 -718 292 -646
rect 388 -718 400 -646
rect 280 -1734 400 -718
rect 280 -1806 292 -1734
rect 388 -1806 400 -1734
rect 280 -2822 400 -1806
rect 280 -2894 292 -2822
rect 388 -2894 400 -2822
rect 280 -2906 400 -2894
rect 2978 -102 3098 454
rect 2978 -174 2990 -102
rect 3086 -174 3098 -102
rect 2978 -1190 3098 -174
rect 2978 -1262 2990 -1190
rect 3086 -1262 3098 -1190
rect 2978 -2278 3098 -1262
rect 2978 -2350 2990 -2278
rect 3086 -2350 3098 -2278
rect 2978 -2906 3098 -2350
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_4 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624298412
transform 1 0 -2242 0 1 -2314
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_5
timestamp 1624298412
transform 1 0 -2242 0 -1 -2314
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624298412
transform 1 0 -2584 0 1 -2314
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1624298412
transform 1 0 -2584 0 -1 -2314
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_9
timestamp 1624298412
transform 1 0 456 0 1 -2314
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_10
timestamp 1624298412
transform 1 0 456 0 -1 -2314
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_5 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624298412
transform 1 0 -218 0 -1 -2314
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_4
timestamp 1624298412
transform 1 0 -218 0 1 -2314
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_5 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624299007
transform 1 0 -494 0 -1 -2314
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_4
timestamp 1624299007
transform 1 0 -494 0 1 -2314
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_10
timestamp 1624298412
transform 1 0 2480 0 -1 -2314
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_9
timestamp 1624298412
transform 1 0 2480 0 1 -2314
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_10
timestamp 1624299007
transform 1 0 2204 0 -1 -2314
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_9
timestamp 1624299007
transform 1 0 2204 0 1 -2314
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1624298412
transform -1 0 3282 0 1 -2314
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1624298412
transform -1 0 3282 0 -1 -2314
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1624298412
transform 1 0 -2242 0 -1 -1226
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1624298412
transform 1 0 -2584 0 -1 -1226
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_8
timestamp 1624298412
transform 1 0 456 0 -1 -1226
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_2
timestamp 1624298412
transform 1 0 -218 0 -1 -1226
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1624299007
transform 1 0 -494 0 -1 -1226
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_8
timestamp 1624298412
transform 1 0 2480 0 -1 -1226
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_8
timestamp 1624299007
transform 1 0 2204 0 -1 -1226
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1624298412
transform -1 0 3282 0 -1 -1226
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1624298412
transform 1 0 -2242 0 1 -1226
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1624298412
transform 1 0 -2584 0 1 -1226
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_7
timestamp 1624298412
transform 1 0 456 0 1 -1226
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_3
timestamp 1624298412
transform 1 0 -218 0 1 -1226
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1624299007
transform 1 0 -494 0 1 -1226
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_7
timestamp 1624298412
transform 1 0 2480 0 1 -1226
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_7
timestamp 1624299007
transform 1 0 2204 0 1 -1226
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1624298412
transform -1 0 3282 0 1 -1226
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1
timestamp 1624298412
transform 1 0 -2242 0 -1 -138
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1624298412
transform 1 0 -2584 0 -1 -138
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_6
timestamp 1624298412
transform 1 0 456 0 -1 -138
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_1
timestamp 1624298412
transform 1 0 -218 0 -1 -138
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1624299007
transform 1 0 -494 0 -1 -138
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_6
timestamp 1624298412
transform 1 0 2480 0 -1 -138
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_6
timestamp 1624299007
transform 1 0 2204 0 -1 -138
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1624298412
transform -1 0 3282 0 -1 -138
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_0
timestamp 1624298412
transform 1 0 -2242 0 1 -138
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1624298412
transform 1 0 -2584 0 1 -138
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  sky130_fd_sc_hd__inv_4_0
timestamp 1624298412
transform 1 0 -218 0 1 -138
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1624298412
transform 1 0 316 0 1 -138
box -38 -48 130 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1624299007
transform 1 0 -494 0 1 -138
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1624298412
transform -1 0 3282 0 1 -138
box -38 -48 130 592
<< labels >>
rlabel comment s -2242 -1226 -2242 -1226 4 dfxbp_1
rlabel comment s -2242 -2314 -2242 -2314 4 dfxbp_1
flabel metal1 s -2562 -691 -2509 -662 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel comment s -2584 -138 -2584 -138 2 tapvpwrvgnd_1
flabel metal1 s -2562 -702 -2509 -673 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s -2562 -1779 -2509 -1750 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel comment s -2584 -1226 -2584 -1226 2 tapvpwrvgnd_1
flabel metal1 s -2562 -1790 -2509 -1761 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s -2562 -2867 -2509 -2838 0 FreeSans 200 0 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel comment s -2584 -2314 -2584 -2314 2 tapvpwrvgnd_1
rlabel comment s 3282 -2314 3282 -2314 8 tapvpwrvgnd_1
flabel metal1 s 3207 -2867 3260 -2838 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 3207 -1790 3260 -1761 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel comment s 3282 -1226 3282 -1226 8 tapvpwrvgnd_1
flabel metal1 s 3207 -1779 3260 -1750 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 s 3207 -702 3260 -673 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
rlabel comment s 3282 -138 3282 -138 8 tapvpwrvgnd_1
flabel metal1 s 3207 -691 3260 -662 0 FreeSans 200 180 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel metal1 -2660 116 -2654 122 1 FreeSans 480 0 0 0 vin
flabel metal1 s 3210 -1244 3261 -1206 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 3210 -1246 3261 -1208 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 3210 -2332 3261 -2294 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 3210 -2334 3261 -2296 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s -2563 -2334 -2512 -2296 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s -2563 -2332 -2512 -2294 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s -2563 -1246 -2512 -1208 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s -2563 -1244 -2512 -1206 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s -2563 -158 -2512 -120 0 FreeSans 200 0 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 3210 -158 3261 -120 0 FreeSans 200 180 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal4 -2348 -374 -2344 -370 1 FreeSans 480 0 0 0 VSS
flabel metal4 332 -378 342 -370 1 FreeSans 480 0 0 0 VDD
flabel metal2 1856 80 1866 88 1 FreeSans 480 0 0 0 vout
<< end >>

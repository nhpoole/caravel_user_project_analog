magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nmos >>
rect -2545 109 -1745 309
rect -1687 109 -887 309
rect -829 109 -29 309
rect 29 109 829 309
rect 887 109 1687 309
rect 1745 109 2545 309
rect -2545 -309 -1745 -109
rect -1687 -309 -887 -109
rect -829 -309 -29 -109
rect 29 -309 829 -109
rect 887 -309 1687 -109
rect 1745 -309 2545 -109
<< ndiff >>
rect -2603 297 -2545 309
rect -2603 121 -2591 297
rect -2557 121 -2545 297
rect -2603 109 -2545 121
rect -1745 297 -1687 309
rect -1745 121 -1733 297
rect -1699 121 -1687 297
rect -1745 109 -1687 121
rect -887 297 -829 309
rect -887 121 -875 297
rect -841 121 -829 297
rect -887 109 -829 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 829 297 887 309
rect 829 121 841 297
rect 875 121 887 297
rect 829 109 887 121
rect 1687 297 1745 309
rect 1687 121 1699 297
rect 1733 121 1745 297
rect 1687 109 1745 121
rect 2545 297 2603 309
rect 2545 121 2557 297
rect 2591 121 2603 297
rect 2545 109 2603 121
rect -2603 -121 -2545 -109
rect -2603 -297 -2591 -121
rect -2557 -297 -2545 -121
rect -2603 -309 -2545 -297
rect -1745 -121 -1687 -109
rect -1745 -297 -1733 -121
rect -1699 -297 -1687 -121
rect -1745 -309 -1687 -297
rect -887 -121 -829 -109
rect -887 -297 -875 -121
rect -841 -297 -829 -121
rect -887 -309 -829 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 829 -121 887 -109
rect 829 -297 841 -121
rect 875 -297 887 -121
rect 829 -309 887 -297
rect 1687 -121 1745 -109
rect 1687 -297 1699 -121
rect 1733 -297 1745 -121
rect 1687 -309 1745 -297
rect 2545 -121 2603 -109
rect 2545 -297 2557 -121
rect 2591 -297 2603 -121
rect 2545 -309 2603 -297
<< ndiffc >>
rect -2591 121 -2557 297
rect -1733 121 -1699 297
rect -875 121 -841 297
rect -17 121 17 297
rect 841 121 875 297
rect 1699 121 1733 297
rect 2557 121 2591 297
rect -2591 -297 -2557 -121
rect -1733 -297 -1699 -121
rect -875 -297 -841 -121
rect -17 -297 17 -121
rect 841 -297 875 -121
rect 1699 -297 1733 -121
rect 2557 -297 2591 -121
<< poly >>
rect -2391 381 -1899 397
rect -2391 364 -2375 381
rect -2545 347 -2375 364
rect -1915 364 -1899 381
rect -1533 381 -1041 397
rect -1533 364 -1517 381
rect -1915 347 -1745 364
rect -2545 309 -1745 347
rect -1687 347 -1517 364
rect -1057 364 -1041 381
rect -675 381 -183 397
rect -675 364 -659 381
rect -1057 347 -887 364
rect -1687 309 -887 347
rect -829 347 -659 364
rect -199 364 -183 381
rect 183 381 675 397
rect 183 364 199 381
rect -199 347 -29 364
rect -829 309 -29 347
rect 29 347 199 364
rect 659 364 675 381
rect 1041 381 1533 397
rect 1041 364 1057 381
rect 659 347 829 364
rect 29 309 829 347
rect 887 347 1057 364
rect 1517 364 1533 381
rect 1899 381 2391 397
rect 1899 364 1915 381
rect 1517 347 1687 364
rect 887 309 1687 347
rect 1745 347 1915 364
rect 2375 364 2391 381
rect 2375 347 2545 364
rect 1745 309 2545 347
rect -2545 71 -1745 109
rect -2545 54 -2375 71
rect -2391 37 -2375 54
rect -1915 54 -1745 71
rect -1687 71 -887 109
rect -1687 54 -1517 71
rect -1915 37 -1899 54
rect -2391 21 -1899 37
rect -1533 37 -1517 54
rect -1057 54 -887 71
rect -829 71 -29 109
rect -829 54 -659 71
rect -1057 37 -1041 54
rect -1533 21 -1041 37
rect -675 37 -659 54
rect -199 54 -29 71
rect 29 71 829 109
rect 29 54 199 71
rect -199 37 -183 54
rect -675 21 -183 37
rect 183 37 199 54
rect 659 54 829 71
rect 887 71 1687 109
rect 887 54 1057 71
rect 659 37 675 54
rect 183 21 675 37
rect 1041 37 1057 54
rect 1517 54 1687 71
rect 1745 71 2545 109
rect 1745 54 1915 71
rect 1517 37 1533 54
rect 1041 21 1533 37
rect 1899 37 1915 54
rect 2375 54 2545 71
rect 2375 37 2391 54
rect 1899 21 2391 37
rect -2391 -37 -1899 -21
rect -2391 -54 -2375 -37
rect -2545 -71 -2375 -54
rect -1915 -54 -1899 -37
rect -1533 -37 -1041 -21
rect -1533 -54 -1517 -37
rect -1915 -71 -1745 -54
rect -2545 -109 -1745 -71
rect -1687 -71 -1517 -54
rect -1057 -54 -1041 -37
rect -675 -37 -183 -21
rect -675 -54 -659 -37
rect -1057 -71 -887 -54
rect -1687 -109 -887 -71
rect -829 -71 -659 -54
rect -199 -54 -183 -37
rect 183 -37 675 -21
rect 183 -54 199 -37
rect -199 -71 -29 -54
rect -829 -109 -29 -71
rect 29 -71 199 -54
rect 659 -54 675 -37
rect 1041 -37 1533 -21
rect 1041 -54 1057 -37
rect 659 -71 829 -54
rect 29 -109 829 -71
rect 887 -71 1057 -54
rect 1517 -54 1533 -37
rect 1899 -37 2391 -21
rect 1899 -54 1915 -37
rect 1517 -71 1687 -54
rect 887 -109 1687 -71
rect 1745 -71 1915 -54
rect 2375 -54 2391 -37
rect 2375 -71 2545 -54
rect 1745 -109 2545 -71
rect -2545 -347 -1745 -309
rect -2545 -364 -2375 -347
rect -2391 -381 -2375 -364
rect -1915 -364 -1745 -347
rect -1687 -347 -887 -309
rect -1687 -364 -1517 -347
rect -1915 -381 -1899 -364
rect -2391 -397 -1899 -381
rect -1533 -381 -1517 -364
rect -1057 -364 -887 -347
rect -829 -347 -29 -309
rect -829 -364 -659 -347
rect -1057 -381 -1041 -364
rect -1533 -397 -1041 -381
rect -675 -381 -659 -364
rect -199 -364 -29 -347
rect 29 -347 829 -309
rect 29 -364 199 -347
rect -199 -381 -183 -364
rect -675 -397 -183 -381
rect 183 -381 199 -364
rect 659 -364 829 -347
rect 887 -347 1687 -309
rect 887 -364 1057 -347
rect 659 -381 675 -364
rect 183 -397 675 -381
rect 1041 -381 1057 -364
rect 1517 -364 1687 -347
rect 1745 -347 2545 -309
rect 1745 -364 1915 -347
rect 1517 -381 1533 -364
rect 1041 -397 1533 -381
rect 1899 -381 1915 -364
rect 2375 -364 2545 -347
rect 2375 -381 2391 -364
rect 1899 -397 2391 -381
<< polycont >>
rect -2375 347 -1915 381
rect -1517 347 -1057 381
rect -659 347 -199 381
rect 199 347 659 381
rect 1057 347 1517 381
rect 1915 347 2375 381
rect -2375 37 -1915 71
rect -1517 37 -1057 71
rect -659 37 -199 71
rect 199 37 659 71
rect 1057 37 1517 71
rect 1915 37 2375 71
rect -2375 -71 -1915 -37
rect -1517 -71 -1057 -37
rect -659 -71 -199 -37
rect 199 -71 659 -37
rect 1057 -71 1517 -37
rect 1915 -71 2375 -37
rect -2375 -381 -1915 -347
rect -1517 -381 -1057 -347
rect -659 -381 -199 -347
rect 199 -381 659 -347
rect 1057 -381 1517 -347
rect 1915 -381 2375 -347
<< locali >>
rect -2391 347 -2375 381
rect -1915 347 -1899 381
rect -1533 347 -1517 381
rect -1057 347 -1041 381
rect -675 347 -659 381
rect -199 347 -183 381
rect 183 347 199 381
rect 659 347 675 381
rect 1041 347 1057 381
rect 1517 347 1533 381
rect 1899 347 1915 381
rect 2375 347 2391 381
rect -2591 297 -2557 313
rect -2591 105 -2557 121
rect -1733 297 -1699 313
rect -1733 105 -1699 121
rect -875 297 -841 313
rect -875 105 -841 121
rect -17 297 17 313
rect -17 105 17 121
rect 841 297 875 313
rect 841 105 875 121
rect 1699 297 1733 313
rect 1699 105 1733 121
rect 2557 297 2591 313
rect 2557 105 2591 121
rect -2391 37 -2375 71
rect -1915 37 -1899 71
rect -1533 37 -1517 71
rect -1057 37 -1041 71
rect -675 37 -659 71
rect -199 37 -183 71
rect 183 37 199 71
rect 659 37 675 71
rect 1041 37 1057 71
rect 1517 37 1533 71
rect 1899 37 1915 71
rect 2375 37 2391 71
rect -2391 -71 -2375 -37
rect -1915 -71 -1899 -37
rect -1533 -71 -1517 -37
rect -1057 -71 -1041 -37
rect -675 -71 -659 -37
rect -199 -71 -183 -37
rect 183 -71 199 -37
rect 659 -71 675 -37
rect 1041 -71 1057 -37
rect 1517 -71 1533 -37
rect 1899 -71 1915 -37
rect 2375 -71 2391 -37
rect -2591 -121 -2557 -105
rect -2591 -313 -2557 -297
rect -1733 -121 -1699 -105
rect -1733 -313 -1699 -297
rect -875 -121 -841 -105
rect -875 -313 -841 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 841 -121 875 -105
rect 841 -313 875 -297
rect 1699 -121 1733 -105
rect 1699 -313 1733 -297
rect 2557 -121 2591 -105
rect 2557 -313 2591 -297
rect -2391 -381 -2375 -347
rect -1915 -381 -1899 -347
rect -1533 -381 -1517 -347
rect -1057 -381 -1041 -347
rect -675 -381 -659 -347
rect -199 -381 -183 -347
rect 183 -381 199 -347
rect 659 -381 675 -347
rect 1041 -381 1057 -347
rect 1517 -381 1533 -347
rect 1899 -381 1915 -347
rect 2375 -381 2391 -347
<< viali >>
rect -2337 347 -1953 381
rect -1479 347 -1095 381
rect -621 347 -237 381
rect 237 347 621 381
rect 1095 347 1479 381
rect 1953 347 2337 381
rect -2591 121 -2557 297
rect -1733 121 -1699 297
rect -875 121 -841 297
rect -17 121 17 297
rect 841 121 875 297
rect 1699 121 1733 297
rect 2557 121 2591 297
rect -2337 37 -1953 71
rect -1479 37 -1095 71
rect -621 37 -237 71
rect 237 37 621 71
rect 1095 37 1479 71
rect 1953 37 2337 71
rect -2337 -71 -1953 -37
rect -1479 -71 -1095 -37
rect -621 -71 -237 -37
rect 237 -71 621 -37
rect 1095 -71 1479 -37
rect 1953 -71 2337 -37
rect -2591 -297 -2557 -121
rect -1733 -297 -1699 -121
rect -875 -297 -841 -121
rect -17 -297 17 -121
rect 841 -297 875 -121
rect 1699 -297 1733 -121
rect 2557 -297 2591 -121
rect -2337 -381 -1953 -347
rect -1479 -381 -1095 -347
rect -621 -381 -237 -347
rect 237 -381 621 -347
rect 1095 -381 1479 -347
rect 1953 -381 2337 -347
<< metal1 >>
rect -2349 381 -1941 387
rect -2349 347 -2337 381
rect -1953 347 -1941 381
rect -2349 341 -1941 347
rect -1491 381 -1083 387
rect -1491 347 -1479 381
rect -1095 347 -1083 381
rect -1491 341 -1083 347
rect -633 381 -225 387
rect -633 347 -621 381
rect -237 347 -225 381
rect -633 341 -225 347
rect 225 381 633 387
rect 225 347 237 381
rect 621 347 633 381
rect 225 341 633 347
rect 1083 381 1491 387
rect 1083 347 1095 381
rect 1479 347 1491 381
rect 1083 341 1491 347
rect 1941 381 2349 387
rect 1941 347 1953 381
rect 2337 347 2349 381
rect 1941 341 2349 347
rect -2597 297 -2551 309
rect -2597 121 -2591 297
rect -2557 121 -2551 297
rect -2597 109 -2551 121
rect -1739 297 -1693 309
rect -1739 121 -1733 297
rect -1699 121 -1693 297
rect -1739 109 -1693 121
rect -881 297 -835 309
rect -881 121 -875 297
rect -841 121 -835 297
rect -881 109 -835 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 835 297 881 309
rect 835 121 841 297
rect 875 121 881 297
rect 835 109 881 121
rect 1693 297 1739 309
rect 1693 121 1699 297
rect 1733 121 1739 297
rect 1693 109 1739 121
rect 2551 297 2597 309
rect 2551 121 2557 297
rect 2591 121 2597 297
rect 2551 109 2597 121
rect -2349 71 -1941 77
rect -2349 37 -2337 71
rect -1953 37 -1941 71
rect -2349 31 -1941 37
rect -1491 71 -1083 77
rect -1491 37 -1479 71
rect -1095 37 -1083 71
rect -1491 31 -1083 37
rect -633 71 -225 77
rect -633 37 -621 71
rect -237 37 -225 71
rect -633 31 -225 37
rect 225 71 633 77
rect 225 37 237 71
rect 621 37 633 71
rect 225 31 633 37
rect 1083 71 1491 77
rect 1083 37 1095 71
rect 1479 37 1491 71
rect 1083 31 1491 37
rect 1941 71 2349 77
rect 1941 37 1953 71
rect 2337 37 2349 71
rect 1941 31 2349 37
rect -2349 -37 -1941 -31
rect -2349 -71 -2337 -37
rect -1953 -71 -1941 -37
rect -2349 -77 -1941 -71
rect -1491 -37 -1083 -31
rect -1491 -71 -1479 -37
rect -1095 -71 -1083 -37
rect -1491 -77 -1083 -71
rect -633 -37 -225 -31
rect -633 -71 -621 -37
rect -237 -71 -225 -37
rect -633 -77 -225 -71
rect 225 -37 633 -31
rect 225 -71 237 -37
rect 621 -71 633 -37
rect 225 -77 633 -71
rect 1083 -37 1491 -31
rect 1083 -71 1095 -37
rect 1479 -71 1491 -37
rect 1083 -77 1491 -71
rect 1941 -37 2349 -31
rect 1941 -71 1953 -37
rect 2337 -71 2349 -37
rect 1941 -77 2349 -71
rect -2597 -121 -2551 -109
rect -2597 -297 -2591 -121
rect -2557 -297 -2551 -121
rect -2597 -309 -2551 -297
rect -1739 -121 -1693 -109
rect -1739 -297 -1733 -121
rect -1699 -297 -1693 -121
rect -1739 -309 -1693 -297
rect -881 -121 -835 -109
rect -881 -297 -875 -121
rect -841 -297 -835 -121
rect -881 -309 -835 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 835 -121 881 -109
rect 835 -297 841 -121
rect 875 -297 881 -121
rect 835 -309 881 -297
rect 1693 -121 1739 -109
rect 1693 -297 1699 -121
rect 1733 -297 1739 -121
rect 1693 -309 1739 -297
rect 2551 -121 2597 -109
rect 2551 -297 2557 -121
rect 2591 -297 2597 -121
rect 2551 -309 2597 -297
rect -2349 -347 -1941 -341
rect -2349 -381 -2337 -347
rect -1953 -381 -1941 -347
rect -2349 -387 -1941 -381
rect -1491 -347 -1083 -341
rect -1491 -381 -1479 -347
rect -1095 -381 -1083 -347
rect -1491 -387 -1083 -381
rect -633 -347 -225 -341
rect -633 -381 -621 -347
rect -237 -381 -225 -347
rect -633 -387 -225 -381
rect 225 -347 633 -341
rect 225 -381 237 -347
rect 621 -381 633 -347
rect 225 -387 633 -381
rect 1083 -347 1491 -341
rect 1083 -381 1095 -347
rect 1479 -381 1491 -347
rect 1083 -387 1491 -381
rect 1941 -347 2349 -341
rect 1941 -381 1953 -347
rect 2337 -381 2349 -347
rect 1941 -387 2349 -381
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 1 l 4 m 2 nf 6 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>

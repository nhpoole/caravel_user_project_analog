magic
tech sky130A
magscale 1 2
timestamp 1624298412
<< pwell >>
rect -238 -2078 4438 978
<< psubdiff >>
rect -202 842 -40 942
rect 4240 842 4402 942
rect -202 780 -102 842
rect -202 -1942 -102 -1880
rect 4302 780 4402 842
rect 4302 -1942 4402 -1880
rect -202 -2042 -40 -1942
rect 4240 -2042 4402 -1942
<< psubdiffcont >>
rect -40 842 4240 942
rect -202 -1880 -102 780
rect 4302 -1880 4402 780
rect -40 -2042 4240 -1942
<< locali >>
rect -202 780 -102 942
rect -202 -2042 -102 -1880
rect 4302 780 4402 942
rect 4302 -2042 4402 -1880
<< viali >>
rect -102 842 -40 942
rect -40 842 4240 942
rect 4240 842 4302 942
rect -202 -1773 -102 673
rect 4302 -1773 4402 673
rect -102 -2042 -40 -1942
rect -40 -2042 4240 -1942
rect 4240 -2042 4302 -1942
<< metal1 >>
rect 4662 12790 5100 12860
rect 4662 1198 4704 12790
rect 4962 1198 5100 12790
rect 4662 1148 5100 1198
rect -210 986 4968 1022
rect -210 896 -156 986
rect 4924 896 4968 986
rect -210 842 -102 896
rect 4302 842 4968 896
rect -210 838 4968 842
rect -208 836 4408 838
rect -208 673 -96 836
rect -8 688 -2 748
rect 58 688 64 748
rect -208 -1773 -202 673
rect -102 -1773 -96 673
rect -2 -1218 58 688
rect 136 564 142 624
rect 202 564 208 624
rect 272 620 332 836
rect 404 620 464 836
rect 784 688 790 748
rect 850 688 856 748
rect 142 -1092 202 564
rect 272 560 464 620
rect 272 -244 332 560
rect 404 478 464 560
rect 790 382 850 688
rect 1172 624 1232 836
rect 1304 624 1364 836
rect 1432 624 1492 836
rect 1172 564 1492 624
rect 1812 564 1818 624
rect 1878 564 1884 624
rect 2332 564 2338 624
rect 2398 564 2404 624
rect 2724 622 2784 836
rect 2856 622 2916 836
rect 2984 622 3044 836
rect 3360 688 3366 748
rect 3426 688 3432 748
rect 1172 480 1232 564
rect 1304 562 1492 564
rect 404 -244 464 6
rect 272 -304 464 -244
rect 272 -1090 332 -304
rect 404 -520 464 -304
rect 532 -358 592 80
rect 662 -110 722 4
rect 920 -108 980 0
rect 656 -170 662 -110
rect 722 -170 728 -110
rect 914 -168 920 -108
rect 980 -168 986 -108
rect 526 -418 532 -358
rect 592 -418 598 -358
rect 662 -520 722 -170
rect 784 -300 790 -240
rect 850 -300 856 -240
rect 790 -620 850 -300
rect 920 -518 980 -168
rect 1050 -358 1110 102
rect 1172 -242 1232 6
rect 1304 -242 1364 562
rect 1432 482 1492 562
rect 1818 386 1878 564
rect 2338 390 2398 564
rect 2724 562 3044 622
rect 2724 478 2784 562
rect 2856 560 3044 562
rect 1172 -244 1364 -242
rect 1434 -244 1494 6
rect 1564 -240 1624 104
rect 1692 -110 1752 2
rect 1952 -110 2012 4
rect 1686 -170 1692 -110
rect 1752 -170 1758 -110
rect 1946 -170 1952 -110
rect 2012 -170 2018 -110
rect 1172 -302 1494 -244
rect 1558 -300 1564 -240
rect 1624 -300 1630 -240
rect 1044 -418 1050 -358
rect 1110 -418 1116 -358
rect 1172 -518 1232 -302
rect 1304 -304 1494 -302
rect 398 -1090 458 -994
rect 136 -1152 142 -1092
rect 202 -1152 208 -1092
rect 272 -1150 458 -1090
rect 532 -1092 592 -902
rect 1048 -1092 1108 -910
rect 1170 -1092 1230 -992
rect 1304 -1092 1364 -304
rect 1434 -516 1494 -304
rect 1692 -522 1752 -170
rect 1816 -418 1822 -358
rect 1882 -418 1888 -358
rect 1822 -616 1882 -418
rect 1952 -522 2012 -170
rect 2080 -240 2140 110
rect 2208 -110 2268 8
rect 2466 -110 2526 10
rect 2202 -170 2208 -110
rect 2268 -170 2274 -110
rect 2460 -170 2466 -110
rect 2526 -170 2532 -110
rect 2074 -300 2080 -240
rect 2140 -300 2146 -240
rect 2208 -522 2268 -170
rect 2330 -418 2336 -358
rect 2396 -418 2402 -358
rect 2336 -616 2396 -418
rect 2466 -522 2526 -170
rect 2598 -240 2658 120
rect 2592 -300 2598 -240
rect 2658 -300 2664 -240
rect 2724 -244 2784 4
rect 2856 -244 2916 560
rect 2984 480 3044 560
rect 3366 370 3426 688
rect 3758 624 3818 836
rect 3882 624 3942 836
rect 4128 688 4134 748
rect 4194 688 4200 748
rect 3758 564 3942 624
rect 3992 564 3998 624
rect 4058 564 4064 624
rect 3758 480 3818 564
rect 2724 -246 2916 -244
rect 2986 -246 3046 4
rect 2724 -304 3046 -246
rect 2724 -520 2784 -304
rect 2856 -306 3046 -304
rect 1432 -1092 1492 -992
rect -8 -1278 -2 -1218
rect 58 -1278 64 -1218
rect 272 -1352 332 -1150
rect 398 -1352 458 -1150
rect 526 -1152 532 -1092
rect 592 -1152 598 -1092
rect 1042 -1152 1048 -1092
rect 1108 -1152 1114 -1092
rect 1170 -1152 1492 -1092
rect 1170 -1352 1230 -1152
rect 1304 -1352 1364 -1152
rect 1432 -1352 1492 -1152
rect 1560 -1218 1620 -888
rect 2082 -1218 2142 -894
rect 2596 -1218 2656 -890
rect 2722 -1094 2782 -994
rect 2856 -1094 2916 -306
rect 2986 -518 3046 -306
rect 3112 -358 3172 126
rect 3242 -110 3302 -2
rect 3502 -110 3562 4
rect 3236 -170 3242 -110
rect 3302 -170 3308 -110
rect 3496 -170 3502 -110
rect 3562 -170 3568 -110
rect 3106 -418 3112 -358
rect 3172 -418 3178 -358
rect 3242 -520 3302 -170
rect 3362 -300 3368 -240
rect 3428 -300 3434 -240
rect 3368 -632 3428 -300
rect 3502 -520 3562 -170
rect 3626 -358 3686 102
rect 3754 -240 3814 4
rect 3882 -240 3942 564
rect 3754 -300 3942 -240
rect 3620 -418 3626 -358
rect 3686 -418 3692 -358
rect 3754 -518 3814 -300
rect 2984 -1094 3044 -994
rect 3112 -1092 3172 -902
rect 3626 -1092 3686 -906
rect 3752 -1092 3812 -992
rect 3882 -1092 3942 -300
rect 3998 -1092 4058 564
rect 2722 -1154 3044 -1094
rect 3106 -1152 3112 -1092
rect 3172 -1152 3178 -1092
rect 3620 -1152 3626 -1092
rect 3686 -1152 3692 -1092
rect 3752 -1152 3942 -1092
rect 3992 -1152 3998 -1092
rect 4058 -1152 4064 -1092
rect 1554 -1278 1560 -1218
rect 1620 -1278 1626 -1218
rect 2076 -1278 2082 -1218
rect 2142 -1278 2148 -1218
rect 2590 -1278 2596 -1218
rect 2656 -1278 2662 -1218
rect 2722 -1352 2782 -1154
rect 2856 -1352 2916 -1154
rect 2984 -1352 3044 -1154
rect 3752 -1352 3812 -1152
rect 3882 -1352 3942 -1152
rect 4134 -1218 4194 688
rect 4296 673 4408 836
rect 4128 -1278 4134 -1218
rect 4194 -1278 4200 -1218
rect 204 -1402 3996 -1352
rect 204 -1506 258 -1402
rect 3950 -1506 3996 -1402
rect 204 -1550 3996 -1506
rect -208 -1936 -96 -1773
rect 504 -1936 514 -1636
rect 3686 -1936 3696 -1636
rect 4296 -1773 4302 673
rect 4402 -1773 4408 673
rect 6942 104 7222 164
rect 4296 -1936 4408 -1773
rect -208 -1942 4408 -1936
rect -208 -2042 -102 -1942
rect 4302 -2042 4408 -1942
rect -208 -2048 4408 -2042
<< via1 >>
rect 4704 1198 4962 12790
rect -156 942 4924 986
rect -156 896 -102 942
rect -102 896 4302 942
rect 4302 896 4924 942
rect -2 688 58 748
rect 142 564 202 624
rect 790 688 850 748
rect 1818 564 1878 624
rect 2338 564 2398 624
rect 3366 688 3426 748
rect 662 -170 722 -110
rect 920 -168 980 -108
rect 532 -418 592 -358
rect 790 -300 850 -240
rect 1692 -170 1752 -110
rect 1952 -170 2012 -110
rect 1564 -300 1624 -240
rect 1050 -418 1110 -358
rect 142 -1152 202 -1092
rect 1822 -418 1882 -358
rect 2208 -170 2268 -110
rect 2466 -170 2526 -110
rect 2080 -300 2140 -240
rect 2336 -418 2396 -358
rect 2598 -300 2658 -240
rect 4134 688 4194 748
rect 3998 564 4058 624
rect -2 -1278 58 -1218
rect 532 -1152 592 -1092
rect 1048 -1152 1108 -1092
rect 3242 -170 3302 -110
rect 3502 -170 3562 -110
rect 3112 -418 3172 -358
rect 3368 -300 3428 -240
rect 3626 -418 3686 -358
rect 3112 -1152 3172 -1092
rect 3626 -1152 3686 -1092
rect 3998 -1152 4058 -1092
rect 1560 -1278 1620 -1218
rect 2082 -1278 2142 -1218
rect 2596 -1278 2656 -1218
rect 4134 -1278 4194 -1218
rect 258 -1506 3950 -1402
rect -96 -1936 504 -1636
rect 3696 -1936 4296 -1636
<< metal2 >>
rect 4216 12972 5348 13072
rect 1875 12090 1965 12094
rect 4216 12090 4316 12972
rect 1870 12085 4316 12090
rect 1870 11995 1875 12085
rect 1965 11995 4316 12085
rect 1870 11990 4316 11995
rect 4636 12790 5024 12860
rect 1875 11986 1965 11990
rect 1574 9681 1676 9686
rect 1570 9589 1579 9681
rect 1671 9589 1680 9681
rect 1574 9539 1676 9589
rect 919 9437 1676 9539
rect 919 9387 1021 9437
rect 919 9276 1021 9285
rect 1286 4681 1390 4686
rect 1282 4587 1291 4681
rect 1385 4587 1394 4681
rect 1286 4532 1390 4587
rect 1286 4428 1746 4532
rect 1642 4366 1746 4428
rect 1642 4253 1746 4262
rect 4636 1198 4704 12790
rect 4962 1198 5024 12790
rect 5248 12784 5348 12972
rect 5248 12675 5348 12684
rect 4636 1148 5024 1198
rect 5564 1602 8252 1662
rect -202 986 4964 1026
rect -202 896 -156 986
rect 4924 896 4964 986
rect -202 846 4964 896
rect -2 748 58 754
rect 790 748 850 754
rect 3366 748 3426 754
rect 4134 748 4194 754
rect 58 688 790 748
rect 850 688 3366 748
rect 3426 688 4134 748
rect -2 682 58 688
rect 790 682 850 688
rect 3366 682 3426 688
rect 4134 682 4194 688
rect 1033 639 1123 648
rect 142 624 202 630
rect 202 564 1033 624
rect 142 558 202 564
rect 1818 624 1878 630
rect 2338 624 2398 630
rect 3998 624 4058 630
rect 5564 624 5624 1602
rect 6398 640 6596 700
rect 6391 634 6508 640
rect 1123 564 1818 624
rect 1878 564 2338 624
rect 2398 564 3998 624
rect 4058 564 5624 624
rect 1818 558 1878 564
rect 2338 558 2398 564
rect 3998 558 4058 564
rect 1033 540 1123 549
rect 662 -110 722 -104
rect 920 -108 980 -102
rect 722 -168 920 -110
rect 1692 -110 1752 -104
rect 1952 -110 2012 -104
rect 2208 -110 2268 -104
rect 2466 -110 2526 -104
rect 3242 -110 3302 -104
rect 3502 -110 3562 -104
rect 980 -168 1692 -110
rect 722 -170 1692 -168
rect 1752 -170 1952 -110
rect 2012 -170 2208 -110
rect 2268 -170 2466 -110
rect 2526 -170 3242 -110
rect 3302 -170 3502 -110
rect 662 -176 722 -170
rect 920 -174 980 -170
rect 1692 -176 1752 -170
rect 1952 -176 2012 -170
rect 2208 -176 2268 -170
rect 2466 -176 2526 -170
rect 3242 -176 3302 -170
rect 3502 -176 3562 -170
rect 790 -240 850 -234
rect 1564 -240 1624 -234
rect 2080 -240 2140 -234
rect 2598 -240 2658 -234
rect 3368 -240 3428 -234
rect 850 -300 1564 -240
rect 1624 -300 2080 -240
rect 2140 -300 2598 -240
rect 2658 -300 3368 -240
rect 3428 -300 5112 -240
rect 5172 -300 5181 -240
rect 790 -306 850 -300
rect 1564 -306 1624 -300
rect 2080 -306 2140 -300
rect 2598 -306 2658 -300
rect 3368 -306 3428 -300
rect 3607 -341 3697 -332
rect 532 -358 592 -352
rect 1050 -358 1110 -352
rect 1822 -358 1882 -352
rect 2336 -358 2396 -352
rect 3112 -358 3172 -352
rect 6448 -358 6508 634
rect 592 -418 1050 -358
rect 1110 -418 1822 -358
rect 1882 -418 2336 -358
rect 2396 -418 3112 -358
rect 3172 -418 3607 -358
rect 3697 -418 6508 -358
rect 532 -424 592 -418
rect 1050 -424 1110 -418
rect 1822 -424 1882 -418
rect 2336 -424 2396 -418
rect 3112 -424 3172 -418
rect 3607 -440 3697 -431
rect 142 -1092 202 -1086
rect 532 -1092 592 -1086
rect 1048 -1092 1108 -1086
rect 3112 -1092 3172 -1086
rect 3626 -1092 3686 -1086
rect 3998 -1092 4058 -1086
rect 202 -1152 532 -1092
rect 592 -1152 1048 -1092
rect 1108 -1152 3112 -1092
rect 3172 -1152 3626 -1092
rect 3686 -1152 3998 -1092
rect 142 -1158 202 -1152
rect 532 -1158 592 -1152
rect 1048 -1158 1108 -1152
rect 3112 -1158 3172 -1152
rect 3626 -1158 3686 -1152
rect 3998 -1158 4058 -1152
rect -2 -1218 58 -1212
rect 1560 -1218 1620 -1212
rect 2082 -1218 2142 -1212
rect 2596 -1218 2656 -1212
rect 4134 -1218 4194 -1212
rect 58 -1278 1560 -1218
rect 1620 -1278 2082 -1218
rect 2142 -1278 2596 -1218
rect 2656 -1278 4134 -1218
rect -2 -1284 58 -1278
rect 1560 -1284 1620 -1278
rect 2082 -1284 2142 -1278
rect 2596 -1284 2656 -1278
rect 4134 -1284 4194 -1278
rect 204 -1402 3996 -1352
rect 204 -1506 258 -1402
rect 3950 -1506 3996 -1402
rect 204 -1550 3996 -1506
rect -96 -1636 504 -1626
rect -96 -1946 504 -1936
rect 3696 -1636 4296 -1626
rect 3696 -1946 4296 -1936
<< via2 >>
rect 1875 11995 1965 12085
rect 1579 9589 1671 9681
rect 919 9285 1021 9387
rect 1291 4587 1385 4681
rect 1642 4262 1746 4366
rect 4704 1198 4962 12790
rect 5248 12684 5348 12784
rect -156 896 4924 986
rect 1033 549 1123 639
rect 5112 -300 5172 -240
rect 3607 -358 3697 -341
rect 3607 -418 3626 -358
rect 3626 -418 3686 -358
rect 3686 -418 3697 -358
rect 3607 -431 3697 -418
rect 258 -1506 3950 -1402
rect -96 -1936 504 -1636
rect 3696 -1936 4296 -1636
<< metal3 >>
rect 1944 13222 5056 13468
rect 1872 12944 5056 13222
rect -1766 12790 5056 12944
rect -1766 12340 4704 12790
rect -1766 11834 -1052 12340
rect 3922 12198 4704 12340
rect 1870 12085 1970 12090
rect -841 12038 -743 12043
rect 1627 12038 1725 12043
rect -844 12037 1726 12038
rect -844 11939 -841 12037
rect -743 11939 1627 12037
rect 1725 11939 1726 12037
rect -844 11938 1726 11939
rect 1870 11995 1875 12085
rect 1965 11995 1970 12085
rect -841 11933 -743 11938
rect 1627 11933 1725 11938
rect 1870 11834 1970 11995
rect -1766 11818 -734 11834
rect -1766 9672 -736 11818
rect 1890 11744 1970 11834
rect 522 9691 634 9912
rect 517 9672 523 9691
rect -1766 9634 523 9672
rect -1766 4336 -1052 9634
rect 517 9581 523 9634
rect 633 9581 639 9691
rect 1574 9681 1676 9812
rect 756 9634 1166 9672
rect 1574 9589 1579 9681
rect 1671 9589 1676 9681
rect 1574 9584 1676 9589
rect 522 9580 634 9581
rect 914 9387 1026 9392
rect 2088 9387 2200 9388
rect 914 9334 919 9387
rect -804 9285 919 9334
rect 1021 9336 1026 9387
rect 1021 9334 1298 9336
rect 2083 9334 2089 9387
rect 1021 9285 1396 9334
rect -804 4876 1396 9285
rect 1992 9277 2089 9334
rect 2199 9334 2205 9387
rect 3928 9334 4704 12198
rect 2199 9277 4704 9334
rect 1992 7200 4704 9277
rect 1734 6802 4704 7200
rect 1992 5096 4704 6802
rect -804 4844 1224 4876
rect 1286 4844 1396 4876
rect 1286 4681 1390 4844
rect 1286 4587 1291 4681
rect 1385 4587 1390 4681
rect 2112 4665 2204 4880
rect 1286 4582 1390 4587
rect 2107 4575 2113 4665
rect 2203 4575 2209 4665
rect 2358 4643 4704 5096
rect 2112 4574 2204 4575
rect 3922 4404 4704 4643
rect -1766 2134 -478 4336
rect 834 4288 840 4380
rect 932 4288 938 4380
rect 1637 4366 1751 4371
rect 840 4180 932 4288
rect 1637 4262 1642 4366
rect 1746 4262 1751 4366
rect 1637 4257 1751 4262
rect 1642 4150 1746 4257
rect -1766 1726 -1052 2134
rect 1291 2030 1389 2035
rect 1290 2029 1796 2030
rect 1290 1931 1291 2029
rect 1389 1931 1697 2029
rect 1795 1931 1801 2029
rect 1290 1930 1796 1931
rect 1291 1925 1389 1930
rect 3928 1810 4704 4404
rect 3922 1726 4704 1810
rect -1766 1198 4704 1726
rect 4962 1198 5056 12790
rect 5243 12784 5353 12789
rect 5243 12779 5248 12784
rect 5348 12779 5353 12784
rect 5243 12673 5353 12679
rect -1766 1126 5056 1198
rect -242 1124 5056 1126
rect -242 986 5054 1124
rect -242 896 -156 986
rect 4924 896 5054 986
rect -242 818 5054 896
rect 1291 644 1389 649
rect 1028 643 1390 644
rect 1028 639 1291 643
rect 1028 549 1033 639
rect 1123 549 1291 639
rect 1028 545 1291 549
rect 1389 545 1390 643
rect 1028 544 1390 545
rect 1291 539 1389 544
rect 5247 -220 5345 -215
rect 5094 -221 5346 -220
rect 5094 -240 5247 -221
rect 5094 -300 5112 -240
rect 5172 -300 5247 -240
rect 5094 -319 5247 -300
rect 5345 -319 5346 -221
rect 5094 -320 5346 -319
rect 5247 -325 5345 -320
rect 4043 -336 4141 -331
rect 3602 -337 4142 -336
rect 3602 -341 4043 -337
rect 3602 -431 3607 -341
rect 3697 -431 4043 -341
rect 3602 -435 4043 -431
rect 4141 -435 4142 -337
rect 3602 -436 4142 -435
rect 4043 -441 4141 -436
rect 204 -1402 3996 -1352
rect 204 -1506 258 -1402
rect 3950 -1506 3996 -1402
rect 204 -1550 3996 -1506
rect -106 -1636 514 -1631
rect -106 -1936 -96 -1636
rect 504 -1936 514 -1636
rect -106 -1941 514 -1936
rect 3686 -1636 4306 -1631
rect 3686 -1936 3696 -1636
rect 4296 -1936 4306 -1636
rect 3686 -1941 4306 -1936
<< via3 >>
rect -841 11939 -743 12037
rect 1627 11939 1725 12037
rect 523 9581 633 9691
rect 2089 9277 2199 9387
rect 2113 4575 2203 4665
rect 840 4288 932 4380
rect 1291 1931 1389 2029
rect 1697 1931 1795 2029
rect 5243 12684 5248 12779
rect 5248 12684 5348 12779
rect 5348 12684 5353 12779
rect 5243 12679 5353 12684
rect 1291 545 1389 643
rect 5247 -319 5345 -221
rect 4043 -435 4141 -337
rect 258 -1506 3950 -1402
rect -96 -1936 504 -1636
rect 3696 -1936 4296 -1636
<< metal4 >>
rect 1944 28680 2742 29480
rect 17174 13068 17274 13680
rect 15670 12968 17274 13068
rect 15670 12784 15770 12968
rect 5246 12780 15770 12784
rect 5242 12779 15770 12780
rect -1744 12706 -1644 12734
rect -1750 12606 1212 12706
rect 1654 12606 4620 12706
rect 5242 12679 5243 12779
rect 5353 12684 15770 12779
rect 5353 12679 5354 12684
rect 5242 12678 5354 12679
rect -1744 10950 -1644 12606
rect 1238 12182 3888 12282
rect -1110 12037 -742 12038
rect -1110 11939 -841 12037
rect -743 11939 -742 12037
rect -1110 11938 -742 11939
rect -1744 10850 -1318 10950
rect -1744 8336 -1644 10850
rect -1110 9134 -1010 11938
rect 1238 11660 1338 12182
rect 884 11560 1338 11660
rect 1626 12037 1726 12038
rect 1626 11939 1627 12037
rect 1725 11939 1726 12037
rect 1626 11086 1726 11939
rect 522 9691 2200 9692
rect 522 9581 523 9691
rect 633 9581 2200 9691
rect 522 9580 2200 9581
rect 2088 9387 2200 9580
rect 2088 9277 2089 9387
rect 2199 9277 2200 9387
rect 2088 9276 2200 9277
rect 3788 9134 3888 12182
rect 4520 10936 4620 12606
rect 4162 10828 4620 10936
rect -1110 9034 -434 9134
rect 3246 9034 3888 9134
rect 4520 8336 4620 10828
rect -1752 8228 -1294 8336
rect 4162 8228 4620 8336
rect -1744 5836 -1644 8228
rect 246 6546 346 7417
rect 2522 6546 2622 7417
rect -1752 5728 -1294 5836
rect 4520 5736 4620 8228
rect -1744 3236 -1644 5728
rect 4162 5628 4620 5736
rect -1108 4782 -358 4882
rect 3020 4786 3891 4886
rect -1752 3128 -1264 3236
rect -1744 1478 -1644 3128
rect -1108 2030 -1008 4782
rect 2112 4665 2204 4666
rect 2112 4575 2113 4665
rect 2203 4575 2204 4665
rect 839 4380 933 4381
rect 2112 4380 2204 4575
rect 839 4288 840 4380
rect 932 4288 2204 4380
rect 839 4287 933 4288
rect 890 2196 1018 2414
rect 890 2096 1590 2196
rect -1108 2029 1390 2030
rect -1108 1931 1291 2029
rect 1389 1931 1390 2029
rect -1108 1930 1390 1931
rect -1744 1378 1206 1478
rect 1290 643 1390 1930
rect 1490 1840 1590 2096
rect 1696 2029 1796 2654
rect 1696 1931 1697 2029
rect 1795 1931 1796 2029
rect 1696 1930 1796 1931
rect 3791 1840 3891 4786
rect 4520 3236 4620 5628
rect 4162 3128 4620 3236
rect 1490 1740 3891 1840
rect 1490 1140 1590 1740
rect 4520 1478 4620 3128
rect 1658 1378 4620 1478
rect 1490 1040 4142 1140
rect 1290 545 1291 643
rect 1389 545 1390 643
rect 1290 544 1390 545
rect 4042 -337 4142 1040
rect 5246 -221 5346 12678
rect 5246 -319 5247 -221
rect 5345 -319 5346 -221
rect 5246 -320 5346 -319
rect 4042 -435 4043 -337
rect 4141 -435 4142 -337
rect 4042 -436 4142 -435
rect -280 -1402 4480 -1320
rect -280 -1506 258 -1402
rect 3950 -1506 4480 -1402
rect -280 -1636 4480 -1506
rect -280 -1936 -96 -1636
rect 504 -1936 3696 -1636
rect 4296 -1936 4480 -1636
rect -280 -2120 4480 -1936
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_7
timestamp 1624298412
transform 1 0 2628 0 1 3234
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_6
timestamp 1624298412
transform 1 0 106 0 1 3234
box -1150 -1100 1050 1100
use sky130_fd_pr__nfet_01v8_USKJ3F  sky130_fd_pr__nfet_01v8_USKJ3F_1
timestamp 1624298412
transform 1 0 2109 0 1 -758
box -1835 -288 1835 288
use sky130_fd_pr__nfet_01v8_USKJ3F  sky130_fd_pr__nfet_01v8_USKJ3F_0
timestamp 1624298412
transform 1 0 2109 0 1 242
box -1835 -288 1835 288
use sky130_fd_pr__cap_mim_m3_1_XQCLDR  sky130_fd_pr__cap_mim_m3_1_XQCLDR_3
timestamp 1624298412
transform -1 0 -1407 0 -1 3106
box -350 -1300 349 1300
use sky130_fd_pr__cap_mim_m3_1_5E2G4H  sky130_fd_pr__cap_mim_m3_1_5E2G4H_3
timestamp 1624298412
transform -1 0 -203 0 -1 1426
box -1550 -300 1549 300
use sky130_fd_pr__cap_mim_m3_1_5E2G4H  sky130_fd_pr__cap_mim_m3_1_5E2G4H_2
timestamp 1624298412
transform 1 0 3068 0 -1 1426
box -1550 -300 1549 300
use sky130_fd_pr__cap_mim_m3_1_XQCLDR  sky130_fd_pr__cap_mim_m3_1_XQCLDR_2
timestamp 1624298412
transform 1 0 4272 0 -1 3106
box -350 -1300 349 1300
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_3
timestamp 1624298412
transform -1 0 -1407 0 1 5756
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_0
timestamp 1624298412
transform -1 0 -1407 0 -1 8250
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_5
timestamp 1624298412
transform 1 0 2884 0 1 5734
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_2
timestamp 1624298412
transform 1 0 2884 0 1 8234
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_3
timestamp 1624298412
transform 1 0 346 0 1 8234
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_4
timestamp 1624298412
transform 1 0 346 0 1 5734
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_1
timestamp 1624298412
transform 1 0 4272 0 -1 8250
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_VQCCU2  sky130_fd_pr__cap_mim_m3_1_VQCCU2_2
timestamp 1624298412
transform 1 0 4272 0 1 5756
box -350 -1100 349 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_1
timestamp 1624298412
transform 1 0 2626 0 1 10734
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_KBZ9JD  sky130_fd_pr__cap_mim_m3_1_KBZ9JD_0
timestamp 1624298412
transform 1 0 116 0 1 10734
box -1150 -1100 1050 1100
use sky130_fd_pr__cap_mim_m3_1_XQCLDR  sky130_fd_pr__cap_mim_m3_1_XQCLDR_1
timestamp 1624298412
transform -1 0 -1407 0 1 10900
box -350 -1300 349 1300
use sky130_fd_pr__cap_mim_m3_1_5E2G4H  sky130_fd_pr__cap_mim_m3_1_5E2G4H_1
timestamp 1624298412
transform -1 0 -203 0 1 12640
box -1550 -300 1549 300
use sky130_fd_pr__cap_mim_m3_1_5E2G4H  sky130_fd_pr__cap_mim_m3_1_5E2G4H_0
timestamp 1624298412
transform 1 0 3068 0 1 12640
box -1550 -300 1549 300
use sky130_fd_pr__cap_mim_m3_1_XQCLDR  sky130_fd_pr__cap_mim_m3_1_XQCLDR_0
timestamp 1624298412
transform 1 0 4272 0 1 10900
box -350 -1300 349 1300
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/se_fold_casc_wide_swing_ota
timestamp 1624298412
transform 1 0 17040 0 1 25080
box -15168 -27258 25000 4400
<< labels >>
flabel metal2 2362 -152 2380 -136 1 FreeSans 480 0 0 0 clk
flabel metal2 2348 -280 2366 -264 1 FreeSans 480 0 0 0 vout
flabel metal1 18 -178 30 -162 1 FreeSans 480 0 0 0 vin
flabel metal2 1848 -1132 1870 -1116 1 FreeSans 480 0 0 0 vholdm
flabel metal2 2620 -404 2638 -386 1 FreeSans 480 0 0 0 vhold
flabel metal4 3836 11340 3852 11354 1 FreeSans 480 0 0 0 vhold
flabel metal1 6974 124 6984 136 1 FreeSans 480 0 0 0 ibiasn
flabel metal4 2134 29128 2186 29174 1 FreeSans 480 0 0 0 VDD
flabel metal4 -1076 11268 -1050 11288 1 FreeSans 480 0 0 0 vholdm
flabel metal3 1324 6968 1358 6998 1 FreeSans 480 0 0 0 vout
flabel metal4 -266 -1346 -260 -1342 1 FreeSans 480 0 0 0 VSS
<< properties >>
string FIXED_BBOX -152 -1992 4352 1492
<< end >>

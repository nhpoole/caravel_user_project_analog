magic
tech sky130A
magscale 1 2
timestamp 1624134973
<< nwell >>
rect -11247 15506 -9306 16346
rect -7803 15507 -7200 15828
<< viali >>
rect -7288 15458 -7240 15506
rect -7184 15462 -7136 15510
<< metal1 >>
rect -4458 30288 -4398 30294
rect -4458 16436 -4398 30228
rect -11018 16376 -9518 16436
rect -8284 16376 -7916 16436
rect -7856 16376 -7850 16436
rect -4464 16376 -4458 16436
rect -4398 16376 -4392 16436
rect -7540 15742 -7332 15838
rect -7490 15506 -7228 15512
rect -7490 15458 -7288 15506
rect -7240 15458 -7228 15506
rect -7490 15452 -7228 15458
rect -7196 15510 -7030 15516
rect -7196 15462 -7184 15510
rect -7136 15462 -7030 15510
rect -7196 15456 -7030 15462
rect -7528 15198 -7326 15294
rect -9694 14740 -9688 14760
rect -11068 14680 -9566 14740
rect -8452 14680 -1320 14740
rect 664 1564 1066 1624
<< via1 >>
rect -4458 30228 -4398 30288
rect -7916 16376 -7856 16436
rect -4458 16376 -4398 16436
<< metal2 >>
rect -4458 30288 -4398 30297
rect -4464 30228 -4458 30288
rect -4398 30228 -4392 30288
rect -4458 30219 -4398 30228
rect -7916 16436 -7856 16442
rect -4458 16436 -4398 16442
rect -7856 16376 -4458 16436
rect -7916 16370 -7856 16376
rect -4458 16370 -4398 16376
rect -13297 15502 -13288 15562
rect -13228 15502 -11530 15562
rect -9675 15502 -9666 15562
rect -9606 15502 -8926 15562
rect -12495 15353 -12486 15413
rect -12426 15353 -11732 15413
rect -9859 15353 -9850 15413
rect -9790 15353 -9164 15413
rect -10082 14806 -7716 14866
rect -13105 14576 -13015 14580
rect -9874 14576 -9774 14585
rect -13110 14571 -9874 14576
rect -13110 14481 -13105 14571
rect -13015 14481 -9874 14571
rect -13110 14476 -9874 14481
rect -9774 14476 -9766 14576
rect -13105 14472 -13015 14476
rect -9874 14467 -9774 14476
rect -13499 14354 -13409 14358
rect -9686 14354 -9586 14363
rect -13504 14349 -9686 14354
rect -13504 14259 -13499 14349
rect -13409 14259 -9686 14349
rect -13504 14254 -9686 14259
rect -13499 14250 -13409 14254
rect -9686 14245 -9586 14254
rect -1851 6458 -1842 6518
rect -1782 6458 480 6518
rect -1566 5556 -1506 5565
rect -1506 5496 2058 5556
rect -1566 5487 -1506 5496
<< via2 >>
rect -4458 30228 -4398 30288
rect -13288 15502 -13228 15562
rect -9666 15502 -9606 15562
rect -12486 15353 -12426 15413
rect -9850 15353 -9790 15413
rect -13105 14481 -13015 14571
rect -9874 14476 -9774 14576
rect -13499 14259 -13409 14349
rect -9686 14254 -9586 14354
rect -1842 6458 -1782 6518
rect -1566 5496 -1506 5556
<< metal3 >>
rect -4486 30293 -4350 30322
rect -4486 30229 -4463 30293
rect -4393 30229 -4350 30293
rect -4486 30228 -4458 30229
rect -4398 30228 -4350 30229
rect -4486 30192 -4350 30228
rect -13310 15562 -13210 15584
rect -13310 15502 -13288 15562
rect -13228 15502 -13210 15562
rect -13504 14349 -13404 14354
rect -13504 14259 -13499 14349
rect -13409 14259 -13404 14349
rect -13504 3637 -13404 14259
rect -13310 5795 -13210 15502
rect -9686 15562 -9586 15580
rect -9686 15502 -9666 15562
rect -9606 15502 -9586 15562
rect -12510 15413 -12410 15434
rect -12510 15353 -12486 15413
rect -12426 15353 -12410 15413
rect -13110 14571 -13010 14576
rect -13110 14481 -13105 14571
rect -13015 14481 -13010 14571
rect -13110 10875 -13010 14481
rect -12510 12903 -12410 15353
rect -9874 15413 -9774 15436
rect -9874 15353 -9850 15413
rect -9790 15353 -9774 15413
rect -9874 14581 -9774 15353
rect -9879 14576 -9769 14581
rect -9879 14476 -9874 14576
rect -9774 14476 -9769 14576
rect -9879 14471 -9769 14476
rect -9686 14359 -9586 15502
rect 10952 14470 11052 14476
rect -1600 14370 10952 14470
rect -9691 14354 -9581 14359
rect -11340 14342 -10740 14348
rect -12325 13742 -11340 13798
rect -9691 14254 -9686 14354
rect -9586 14254 -9581 14354
rect -9691 14249 -9581 14254
rect -8560 14342 -7960 14348
rect -10740 13742 -8560 13798
rect -6972 14344 -6372 14350
rect -7736 13798 -6972 13800
rect -7960 13744 -6972 13798
rect -4192 14344 -3592 14350
rect -6372 13744 -4192 13800
rect -3592 13744 -2607 13800
rect -7960 13742 -2607 13744
rect -12325 13200 -2607 13742
rect -12325 13198 -7666 13200
rect -12515 12805 -12509 12903
rect -12411 12805 -12405 12903
rect -12510 12804 -12410 12805
rect -12325 12164 -11725 13198
rect -12912 11564 -12906 12164
rect -12306 11564 -11725 12164
rect -13115 10777 -13109 10875
rect -13011 10777 -13005 10875
rect -13110 10776 -13010 10777
rect -12325 10086 -11725 11564
rect -9964 12934 -7214 13034
rect -9964 10878 -9864 12934
rect -7314 12716 -7214 12934
rect -3207 12166 -2607 13200
rect -1858 12903 -1758 12904
rect -1863 12805 -1857 12903
rect -1759 12805 -1753 12903
rect -3207 11566 -2626 12166
rect -2026 11566 -2020 12166
rect -10156 10875 -10056 10876
rect -10161 10777 -10155 10875
rect -10057 10777 -10051 10875
rect -9964 10778 -9390 10878
rect -9262 10876 -9162 11114
rect -8101 10882 -8003 10887
rect -7570 10882 -7470 10888
rect -8102 10881 -7570 10882
rect -10156 10588 -10056 10777
rect -10156 10476 -10002 10588
rect -9490 10492 -9390 10778
rect -9268 10776 -9262 10876
rect -9162 10776 -9156 10876
rect -8102 10783 -8101 10881
rect -8003 10783 -7570 10881
rect -8102 10782 -7570 10783
rect -5764 10878 -5664 11128
rect -5956 10875 -5856 10876
rect -8101 10777 -8003 10782
rect -7570 10776 -7470 10782
rect -5961 10777 -5955 10875
rect -5857 10777 -5851 10875
rect -5764 10778 -5190 10878
rect -5062 10876 -4962 11114
rect -3901 10880 -3803 10885
rect -3370 10880 -3270 10886
rect -3902 10879 -3370 10880
rect -7192 10492 -7190 10684
rect -5956 10476 -5856 10777
rect -5290 10684 -5190 10778
rect -5068 10776 -5062 10876
rect -4962 10776 -4956 10876
rect -3902 10781 -3901 10879
rect -3803 10781 -3370 10879
rect -3902 10780 -3370 10781
rect -3901 10775 -3803 10780
rect -3370 10774 -3270 10780
rect -5290 10492 -5192 10684
rect -12922 9486 -12916 10086
rect -12316 9486 -11725 10086
rect -13100 8711 -13000 8712
rect -13105 8613 -13099 8711
rect -13001 8613 -12995 8711
rect -13315 5697 -13309 5795
rect -13211 5697 -13205 5795
rect -13310 5696 -13210 5697
rect -13509 3539 -13503 3637
rect -13405 3539 -13399 3637
rect -13504 3538 -13404 3539
rect -13100 1627 -13000 8613
rect -12325 8460 -11725 9486
rect -10102 8712 -10002 10476
rect -3207 10088 -2607 11566
rect -3207 9488 -2616 10088
rect -2016 9488 -2010 10088
rect -7192 8712 -7092 9154
rect -10510 8612 -10504 8712
rect -10404 8612 -7092 8712
rect -6953 8462 -6351 8464
rect -4183 8462 -3581 8464
rect -3207 8462 -2607 9488
rect -11351 8460 -10749 8462
rect -8581 8460 -7979 8462
rect -7510 8460 -2607 8462
rect -12325 7873 -2607 8460
rect -12325 7871 -4183 7873
rect -12325 7860 -11351 7871
rect -10749 7862 -4183 7871
rect -10749 7860 -6351 7862
rect -11351 7263 -10749 7269
rect -8581 7851 -7979 7860
rect -8581 7243 -7979 7249
rect -6953 7853 -6351 7860
rect -6351 7251 -6332 7538
rect -3581 7862 -2607 7873
rect -4183 7265 -3581 7271
rect -6953 7245 -6332 7251
rect -6932 7112 -6332 7245
rect -11324 7104 -10724 7110
rect -12309 6504 -11324 6560
rect -8544 7104 -7944 7110
rect -10724 6504 -8544 6560
rect -6956 7106 -6332 7112
rect -7720 6560 -6956 6562
rect -7944 6506 -6956 6560
rect -6356 6562 -6332 7106
rect -4176 7106 -3576 7112
rect -6356 6506 -4176 6562
rect -3576 6506 -2591 6562
rect -7944 6504 -2591 6506
rect -12309 5962 -2591 6504
rect -12309 5960 -7650 5962
rect -12309 4926 -11709 5960
rect -11490 5696 -11484 5796
rect -11384 5696 -7198 5796
rect -12896 4326 -12890 4926
rect -12290 4326 -11709 4926
rect -12309 2848 -11709 4326
rect -9948 3640 -9848 5696
rect -7298 5478 -7198 5696
rect -3191 4928 -2591 5962
rect -1858 6518 -1758 12805
rect -1600 8863 -1500 14370
rect 10952 14364 11052 14370
rect -1605 8765 -1599 8863
rect -1501 8765 -1495 8863
rect -1600 8764 -1500 8765
rect -1858 6458 -1842 6518
rect -1782 6458 -1758 6518
rect -1858 5665 -1758 6458
rect -1863 5567 -1857 5665
rect -1759 5567 -1753 5665
rect -1858 5566 -1758 5567
rect -1586 5556 -1486 5594
rect -1586 5496 -1566 5556
rect -1506 5496 -1486 5556
rect -3191 4328 -2610 4928
rect -2010 4328 -2004 4928
rect -10140 3637 -10040 3638
rect -10145 3539 -10139 3637
rect -10041 3539 -10035 3637
rect -9948 3540 -9374 3640
rect -9246 3638 -9146 3876
rect -8085 3644 -7987 3649
rect -7554 3644 -7454 3650
rect -8086 3643 -7554 3644
rect -10140 3350 -10040 3539
rect -10140 3238 -9986 3350
rect -9474 3254 -9374 3540
rect -9252 3538 -9246 3638
rect -9146 3538 -9140 3638
rect -8086 3545 -8085 3643
rect -7987 3545 -7554 3643
rect -8086 3544 -7554 3545
rect -5748 3640 -5648 3890
rect -5940 3637 -5840 3638
rect -8085 3539 -7987 3544
rect -7554 3538 -7454 3544
rect -5945 3539 -5939 3637
rect -5841 3539 -5835 3637
rect -5748 3540 -5174 3640
rect -5046 3638 -4946 3876
rect -3885 3644 -3787 3649
rect -3354 3644 -3254 3650
rect -3886 3643 -3354 3644
rect -7176 3254 -7174 3446
rect -5940 3238 -5840 3539
rect -5274 3446 -5174 3540
rect -5052 3538 -5046 3638
rect -4946 3538 -4940 3638
rect -3886 3545 -3885 3643
rect -3787 3545 -3354 3643
rect -3886 3544 -3354 3545
rect -3885 3539 -3787 3544
rect -3354 3538 -3254 3544
rect -5274 3254 -5176 3446
rect -12906 2248 -12900 2848
rect -12300 2248 -11709 2848
rect -13103 1529 -13097 1627
rect -12999 1529 -12993 1627
rect -13100 1528 -13000 1529
rect -12309 1222 -11709 2248
rect -10086 1474 -9986 3238
rect -3191 2850 -2591 4328
rect -3191 2250 -2600 2850
rect -2000 2250 -1994 2850
rect -7176 1474 -7076 1916
rect -10086 1374 -7076 1474
rect -6937 1224 -6335 1226
rect -4167 1224 -3565 1226
rect -3191 1224 -2591 2250
rect -1586 1625 -1486 5496
rect -1591 1527 -1585 1625
rect -1487 1527 -1481 1625
rect -1586 1526 -1486 1527
rect -11335 1222 -10733 1224
rect -8565 1222 -7963 1224
rect -7494 1222 -2591 1224
rect -12309 635 -2591 1222
rect -12309 633 -4167 635
rect -12309 622 -11335 633
rect -10733 624 -4167 633
rect -10733 622 -6335 624
rect -11335 25 -10733 31
rect -8565 613 -7963 622
rect -8565 5 -7963 11
rect -6937 615 -6335 622
rect -3565 624 -2591 635
rect -4167 27 -3565 33
rect -6937 7 -6335 13
<< via3 >>
rect -4463 30288 -4393 30293
rect -4463 30229 -4458 30288
rect -4458 30229 -4398 30288
rect -4398 30229 -4393 30288
rect 10952 14370 11052 14470
rect -11340 13742 -10740 14342
rect -8560 13742 -7960 14342
rect -6972 13744 -6372 14344
rect -4192 13744 -3592 14344
rect -12509 12805 -12411 12903
rect -12906 11564 -12306 12164
rect -13109 10777 -13011 10875
rect -1857 12805 -1759 12903
rect -2626 11566 -2026 12166
rect -10155 10777 -10057 10875
rect -9262 10776 -9162 10876
rect -8101 10783 -8003 10881
rect -7570 10782 -7470 10882
rect -5955 10777 -5857 10875
rect -5062 10776 -4962 10876
rect -3901 10781 -3803 10879
rect -3370 10780 -3270 10880
rect -12916 9486 -12316 10086
rect -13099 8613 -13001 8711
rect -13309 5697 -13211 5795
rect -13503 3539 -13405 3637
rect -2616 9488 -2016 10088
rect -10504 8612 -10404 8712
rect -11351 7269 -10749 7871
rect -8581 7249 -7979 7851
rect -6953 7251 -6351 7853
rect -4183 7271 -3581 7873
rect -11324 6504 -10724 7104
rect -8544 6504 -7944 7104
rect -6956 6506 -6356 7106
rect -4176 6506 -3576 7106
rect -11484 5696 -11384 5796
rect -12890 4326 -12290 4926
rect -1599 8765 -1501 8863
rect -1857 5567 -1759 5665
rect -2610 4328 -2010 4928
rect -10139 3539 -10041 3637
rect -9246 3538 -9146 3638
rect -8085 3545 -7987 3643
rect -7554 3544 -7454 3644
rect -5939 3539 -5841 3637
rect -5046 3538 -4946 3638
rect -3885 3545 -3787 3643
rect -3354 3544 -3254 3644
rect -12900 2248 -12300 2848
rect -13097 1529 -12999 1627
rect -2600 2250 -2000 2850
rect -1585 1527 -1487 1625
rect -11335 31 -10733 633
rect -8565 11 -7963 613
rect -6937 13 -6335 615
rect -4167 33 -3565 635
<< metal4 >>
rect -4928 30293 -3252 30940
rect -4928 30229 -4463 30293
rect -4393 30229 -3252 30293
rect -4928 30140 -3252 30229
rect 10952 14471 11052 15600
rect 10951 14470 11053 14471
rect 10951 14370 10952 14470
rect 11052 14370 11053 14470
rect 10951 14369 11053 14370
rect -6973 14344 -6371 14345
rect -11341 14342 -10739 14343
rect -11341 13742 -11340 14342
rect -10740 13742 -10739 14342
rect -11341 13741 -10739 13742
rect -8561 14342 -7959 14343
rect -8561 13742 -8560 14342
rect -7960 13742 -7959 14342
rect -6973 13744 -6972 14344
rect -6372 13744 -6371 14344
rect -6973 13743 -6371 13744
rect -4193 14344 -3591 14345
rect -4193 13744 -4192 14344
rect -3592 13744 -3591 14344
rect -4193 13743 -3591 13744
rect -8561 13741 -7959 13742
rect -11340 13190 -10740 13741
rect -8560 13180 -7960 13741
rect -6972 13182 -6372 13743
rect -4192 13192 -3592 13743
rect -12510 12903 -1758 12904
rect -12510 12805 -12509 12903
rect -12411 12805 -1857 12903
rect -1759 12805 -1758 12903
rect -12510 12804 -1758 12805
rect -10134 12450 -10034 12804
rect -12907 12164 -12305 12165
rect -12907 11564 -12906 12164
rect -12306 11564 -11734 12164
rect -8246 11784 -7706 11884
rect -12907 11563 -12305 11564
rect -8102 10881 -8002 10882
rect -9263 10876 -9161 10877
rect -13110 10875 -9262 10876
rect -13110 10777 -13109 10875
rect -13011 10777 -10155 10875
rect -10057 10777 -9262 10875
rect -13110 10776 -9262 10777
rect -9162 10776 -9161 10876
rect -9263 10775 -9161 10776
rect -8102 10783 -8101 10881
rect -8003 10783 -8002 10881
rect -8102 10382 -8002 10783
rect -12917 10086 -12315 10087
rect -12917 9486 -12916 10086
rect -12316 9486 -11744 10086
rect -12917 9485 -12315 9486
rect -10152 8864 -10052 9244
rect -7806 8864 -7706 11784
rect -7570 10883 -7470 12804
rect -5934 12450 -5834 12804
rect -4046 11784 -3506 11884
rect -7571 10882 -7469 10883
rect -7571 10782 -7570 10882
rect -7470 10782 -7469 10882
rect -3902 10879 -3802 10880
rect -5063 10876 -4961 10877
rect -7571 10781 -7469 10782
rect -5956 10875 -5062 10876
rect -5956 10777 -5955 10875
rect -5857 10777 -5062 10875
rect -5956 10776 -5062 10777
rect -4962 10776 -4961 10876
rect -5063 10775 -4961 10776
rect -3902 10781 -3901 10879
rect -3803 10781 -3802 10879
rect -3902 10382 -3802 10781
rect -5952 8864 -5852 9244
rect -3606 8864 -3506 11784
rect -3370 10881 -3270 12804
rect -2627 12166 -2025 12167
rect -3198 11566 -2626 12166
rect -2026 11566 -2025 12166
rect -2627 11565 -2025 11566
rect -3371 10880 -3269 10881
rect -3371 10780 -3370 10880
rect -3270 10780 -3269 10880
rect -3371 10779 -3269 10780
rect -2617 10088 -2015 10089
rect -3188 9488 -2616 10088
rect -2016 9488 -2015 10088
rect -2617 9487 -2015 9488
rect -10152 8863 -1500 8864
rect -10152 8765 -1599 8863
rect -1501 8765 -1500 8863
rect -10152 8764 -1500 8765
rect -10505 8712 -10403 8713
rect -13100 8711 -10504 8712
rect -13100 8613 -13099 8711
rect -13001 8613 -10504 8711
rect -13100 8612 -10504 8613
rect -10404 8612 -10403 8712
rect -10505 8611 -10403 8612
rect -11351 7872 -10749 8453
rect -11352 7871 -10748 7872
rect -11352 7269 -11351 7871
rect -10749 7269 -10748 7871
rect -8581 7852 -7979 8423
rect -6953 7854 -6351 8425
rect -4183 7874 -3581 8455
rect -4184 7873 -3580 7874
rect -6954 7853 -6350 7854
rect -11352 7268 -10748 7269
rect -8582 7851 -7978 7852
rect -11306 7105 -10754 7268
rect -8582 7249 -8581 7851
rect -7979 7519 -7978 7851
rect -7979 7249 -7955 7519
rect -6954 7517 -6953 7853
rect -8582 7248 -7955 7249
rect -8517 7105 -7955 7248
rect -6956 7251 -6953 7517
rect -6351 7251 -6350 7853
rect -4184 7271 -4183 7873
rect -3581 7498 -3580 7873
rect -3581 7271 -3576 7498
rect -4184 7270 -3576 7271
rect -6956 7250 -6350 7251
rect -6956 7107 -6394 7250
rect -4128 7107 -3576 7270
rect -6957 7106 -6355 7107
rect -11325 7104 -10723 7105
rect -11325 6504 -11324 7104
rect -10724 6504 -10723 7104
rect -11325 6503 -10723 6504
rect -8545 7104 -7943 7105
rect -8545 6504 -8544 7104
rect -7944 6504 -7943 7104
rect -6957 6506 -6956 7106
rect -6356 6506 -6355 7106
rect -6957 6505 -6355 6506
rect -4177 7106 -3575 7107
rect -4177 6506 -4176 7106
rect -3576 6506 -3575 7106
rect -4177 6505 -3575 6506
rect -8545 6503 -7943 6504
rect -11324 5952 -10724 6503
rect -8544 5942 -7944 6503
rect -6956 5944 -6356 6505
rect -4176 5954 -3576 6505
rect -11485 5796 -11383 5797
rect -13310 5795 -11484 5796
rect -13310 5697 -13309 5795
rect -13211 5697 -11484 5795
rect -13310 5696 -11484 5697
rect -11384 5696 -11383 5796
rect -11485 5695 -11383 5696
rect -10118 5665 -1758 5666
rect -10118 5567 -1857 5665
rect -1759 5567 -1758 5665
rect -10118 5566 -1758 5567
rect -10118 5212 -10018 5566
rect -12891 4926 -12289 4927
rect -12891 4326 -12890 4926
rect -12290 4326 -11718 4926
rect -8230 4546 -7690 4646
rect -12891 4325 -12289 4326
rect -8086 3643 -7986 3644
rect -9247 3638 -9145 3639
rect -13504 3637 -9246 3638
rect -13504 3539 -13503 3637
rect -13405 3539 -10139 3637
rect -10041 3539 -9246 3637
rect -13504 3538 -9246 3539
rect -9146 3538 -9145 3638
rect -9247 3537 -9145 3538
rect -8086 3545 -8085 3643
rect -7987 3545 -7986 3643
rect -8086 3144 -7986 3545
rect -12901 2848 -12299 2849
rect -12901 2248 -12900 2848
rect -12300 2248 -11728 2848
rect -12901 2247 -12299 2248
rect -10136 1628 -10036 2006
rect -13098 1627 -9512 1628
rect -13098 1529 -13097 1627
rect -12999 1626 -9512 1627
rect -7790 1626 -7690 4546
rect -7554 3645 -7454 5566
rect -5918 5212 -5818 5566
rect -4030 4546 -3490 4646
rect -7555 3644 -7453 3645
rect -7555 3544 -7554 3644
rect -7454 3544 -7453 3644
rect -3886 3643 -3786 3644
rect -5047 3638 -4945 3639
rect -7555 3543 -7453 3544
rect -5940 3637 -5046 3638
rect -5940 3539 -5939 3637
rect -5841 3539 -5046 3637
rect -5940 3538 -5046 3539
rect -4946 3538 -4945 3638
rect -5047 3537 -4945 3538
rect -3886 3545 -3885 3643
rect -3787 3545 -3786 3643
rect -3886 3144 -3786 3545
rect -5936 1626 -5836 2006
rect -3590 1626 -3490 4546
rect -3354 3645 -3254 5566
rect -2611 4928 -2009 4929
rect -3182 4328 -2610 4928
rect -2010 4328 -2009 4928
rect -2611 4327 -2009 4328
rect -3355 3644 -3253 3645
rect -3355 3544 -3354 3644
rect -3254 3544 -3253 3644
rect -3355 3543 -3253 3544
rect -2601 2850 -1999 2851
rect -3172 2250 -2600 2850
rect -2000 2250 -1999 2850
rect -2601 2249 -1999 2250
rect -12999 1625 -1486 1626
rect -12999 1529 -1585 1625
rect -13098 1528 -1585 1529
rect -10136 1527 -1585 1528
rect -1487 1527 -1486 1625
rect -10136 1526 -1486 1527
rect -11350 633 -10550 1226
rect -11350 31 -11335 633
rect -10733 140 -10550 633
rect -8608 613 -7937 1231
rect -8608 140 -8565 613
rect -10733 31 -8565 140
rect -11350 11 -8565 31
rect -7963 140 -7937 613
rect -6990 615 -6317 1232
rect -6990 140 -6937 615
rect -7963 13 -6937 140
rect -6335 140 -6317 615
rect -4211 635 -3518 1252
rect -4211 140 -4167 635
rect -6335 33 -4167 140
rect -3565 140 -3518 635
rect -3565 33 -1808 140
rect -6335 13 -1808 33
rect -7963 11 -1808 13
rect -11350 -660 -1808 11
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_0
timestamp 1624127230
transform 1 0 -8594 0 1 924
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_6
timestamp 1624127230
transform 1 0 -10632 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_7
timestamp 1624127230
transform 1 0 -8632 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_4
timestamp 1624127230
transform -1 0 -11077 0 1 924
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_4
timestamp 1624127230
transform 1 0 -11958 0 1 2542
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_8
timestamp 1624127230
transform 1 0 -4432 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_7
timestamp 1624127230
transform 1 0 -3823 0 1 926
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_3
timestamp 1624127230
transform -1 0 -6306 0 1 926
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_9
timestamp 1624127230
transform 1 0 -6432 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_7
timestamp 1624127230
transform -1 0 -2942 0 1 2544
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_5
timestamp 1624127230
transform 1 0 -10632 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_5
timestamp 1624127230
transform 1 0 -11958 0 1 4646
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_4
timestamp 1624127230
transform 1 0 -8632 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_5
timestamp 1624127230
transform -1 0 -11077 0 1 6260
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_1
timestamp 1624127230
transform 1 0 -8594 0 1 6260
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_11
timestamp 1624127230
transform 1 0 -4432 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_10
timestamp 1624127230
transform 1 0 -6432 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_6
timestamp 1624127230
transform 1 0 -3823 0 1 6262
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_2
timestamp 1624127230
transform -1 0 -6306 0 1 6262
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_6
timestamp 1624127230
transform -1 0 -2942 0 1 4648
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_22
timestamp 1624127230
transform 1 0 -11974 0 1 9780
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_46
timestamp 1624127230
transform 1 0 -10648 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_42
timestamp 1624127230
transform 1 0 -8648 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_23
timestamp 1624127230
transform 1 0 -11974 0 1 11884
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_47
timestamp 1624127230
transform 1 0 -10648 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_44
timestamp 1624127230
transform 1 0 -8648 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_23
timestamp 1624127230
transform -1 0 -11093 0 1 8162
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_22
timestamp 1624127230
transform 1 0 -8610 0 1 8162
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_43
timestamp 1624127230
transform 1 0 -6448 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_40
timestamp 1624127230
transform 1 0 -4448 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_45
timestamp 1624127230
transform 1 0 -6448 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_41
timestamp 1624127230
transform 1 0 -4448 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_23
timestamp 1624127230
transform -1 0 -6322 0 1 8164
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_22
timestamp 1624127230
transform 1 0 -3839 0 1 8164
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_20
timestamp 1624127230
transform -1 0 -2958 0 1 9782
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_21
timestamp 1624127230
transform -1 0 -2958 0 1 11886
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_21
timestamp 1624127230
transform -1 0 -11093 0 1 13498
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_20
timestamp 1624127230
transform 1 0 -8610 0 1 13498
box -950 -300 818 300
use txgate  txgate_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/txgate
timestamp 1624127230
transform 1 0 -86501 0 1 -42680
box 74185 57360 76542 59116
use txgate  txgate_1
timestamp 1624127230
transform 1 0 -83901 0 1 -42680
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_21
timestamp 1624127230
transform -1 0 -6322 0 1 13500
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_20
timestamp 1624127230
transform 1 0 -3839 0 1 13500
box -1350 -300 1232 300
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624127230
transform -1 0 -7070 0 1 15246
box -38 -48 314 592
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/se_fold_casc_wide_swing_ota
timestamp 1624132412
transform 1 0 10912 0 1 26540
box -15168 -27258 25000 4400
<< labels >>
flabel metal4 -5616 -342 -5562 -296 1 FreeSans 480 0 0 0 VSS
flabel metal3 -9542 5744 -9520 5764 1 FreeSans 480 0 0 0 vdiffp
flabel metal4 -9662 5600 -9640 5618 1 FreeSans 480 0 0 0 vip
flabel metal4 -9746 1568 -9730 1582 1 FreeSans 480 0 0 0 vim
flabel metal3 -9772 1414 -9760 1428 1 FreeSans 480 0 0 0 vdiffm
flabel metal3 -9862 8658 -9854 8674 1 FreeSans 480 0 0 0 vim
flabel metal4 -9816 8794 -9798 8822 1 FreeSans 480 0 0 0 vse
flabel metal4 -9746 12834 -9732 12846 1 FreeSans 480 0 0 0 vip
flabel metal3 -9752 12980 -9732 12996 1 FreeSans 480 0 0 0 vocm
flabel metal1 704 1582 716 1600 1 FreeSans 480 0 0 0 ibiasn
flabel metal4 -4738 30526 -4712 30558 1 FreeSans 480 0 0 0 VDD
flabel metal1 -7056 15480 -7054 15484 1 FreeSans 480 0 0 0 rst_n
flabel metal1 -7332 15474 -7328 15480 1 FreeSans 480 0 0 0 rst
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< metal3 >>
rect -850 636 849 800
rect -850 -646 765 636
rect 829 -646 849 636
rect -850 -800 849 -646
<< via3 >>
rect 765 -646 829 636
<< mimcap >>
rect -750 660 650 700
rect -750 -660 -710 660
rect 610 -660 650 660
rect -750 -700 650 -660
<< mimcapcontact >>
rect -710 -660 610 660
<< metal4 >>
rect -711 660 611 661
rect -711 -660 -710 660
rect 610 -660 611 660
rect -711 -661 611 -660
rect 749 636 845 662
rect 749 -646 765 636
rect 829 -646 845 636
rect 749 -662 845 -646
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -850 -800 750 800
string parameters w 7.00 l 7.00 val 103.32 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
string library sky130
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nmos >>
rect -3832 -100 -3032 100
rect -2974 -100 -2174 100
rect -2116 -100 -1316 100
rect -1258 -100 -458 100
rect -400 -100 400 100
rect 458 -100 1258 100
rect 1316 -100 2116 100
rect 2174 -100 2974 100
rect 3032 -100 3832 100
<< ndiff >>
rect -3890 88 -3832 100
rect -3890 -88 -3878 88
rect -3844 -88 -3832 88
rect -3890 -100 -3832 -88
rect -3032 88 -2974 100
rect -3032 -88 -3020 88
rect -2986 -88 -2974 88
rect -3032 -100 -2974 -88
rect -2174 88 -2116 100
rect -2174 -88 -2162 88
rect -2128 -88 -2116 88
rect -2174 -100 -2116 -88
rect -1316 88 -1258 100
rect -1316 -88 -1304 88
rect -1270 -88 -1258 88
rect -1316 -100 -1258 -88
rect -458 88 -400 100
rect -458 -88 -446 88
rect -412 -88 -400 88
rect -458 -100 -400 -88
rect 400 88 458 100
rect 400 -88 412 88
rect 446 -88 458 88
rect 400 -100 458 -88
rect 1258 88 1316 100
rect 1258 -88 1270 88
rect 1304 -88 1316 88
rect 1258 -100 1316 -88
rect 2116 88 2174 100
rect 2116 -88 2128 88
rect 2162 -88 2174 88
rect 2116 -100 2174 -88
rect 2974 88 3032 100
rect 2974 -88 2986 88
rect 3020 -88 3032 88
rect 2974 -100 3032 -88
rect 3832 88 3890 100
rect 3832 -88 3844 88
rect 3878 -88 3890 88
rect 3832 -100 3890 -88
<< ndiffc >>
rect -3878 -88 -3844 88
rect -3020 -88 -2986 88
rect -2162 -88 -2128 88
rect -1304 -88 -1270 88
rect -446 -88 -412 88
rect 412 -88 446 88
rect 1270 -88 1304 88
rect 2128 -88 2162 88
rect 2986 -88 3020 88
rect 3844 -88 3878 88
<< poly >>
rect -3678 172 -3186 188
rect -3678 155 -3662 172
rect -3832 138 -3662 155
rect -3202 155 -3186 172
rect -2820 172 -2328 188
rect -2820 155 -2804 172
rect -3202 138 -3032 155
rect -3832 100 -3032 138
rect -2974 138 -2804 155
rect -2344 155 -2328 172
rect -1962 172 -1470 188
rect -1962 155 -1946 172
rect -2344 138 -2174 155
rect -2974 100 -2174 138
rect -2116 138 -1946 155
rect -1486 155 -1470 172
rect -1104 172 -612 188
rect -1104 155 -1088 172
rect -1486 138 -1316 155
rect -2116 100 -1316 138
rect -1258 138 -1088 155
rect -628 155 -612 172
rect -246 172 246 188
rect -246 155 -230 172
rect -628 138 -458 155
rect -1258 100 -458 138
rect -400 138 -230 155
rect 230 155 246 172
rect 612 172 1104 188
rect 612 155 628 172
rect 230 138 400 155
rect -400 100 400 138
rect 458 138 628 155
rect 1088 155 1104 172
rect 1470 172 1962 188
rect 1470 155 1486 172
rect 1088 138 1258 155
rect 458 100 1258 138
rect 1316 138 1486 155
rect 1946 155 1962 172
rect 2328 172 2820 188
rect 2328 155 2344 172
rect 1946 138 2116 155
rect 1316 100 2116 138
rect 2174 138 2344 155
rect 2804 155 2820 172
rect 3186 172 3678 188
rect 3186 155 3202 172
rect 2804 138 2974 155
rect 2174 100 2974 138
rect 3032 138 3202 155
rect 3662 155 3678 172
rect 3662 138 3832 155
rect 3032 100 3832 138
rect -3832 -138 -3032 -100
rect -3832 -155 -3662 -138
rect -3678 -172 -3662 -155
rect -3202 -155 -3032 -138
rect -2974 -138 -2174 -100
rect -2974 -155 -2804 -138
rect -3202 -172 -3186 -155
rect -3678 -188 -3186 -172
rect -2820 -172 -2804 -155
rect -2344 -155 -2174 -138
rect -2116 -138 -1316 -100
rect -2116 -155 -1946 -138
rect -2344 -172 -2328 -155
rect -2820 -188 -2328 -172
rect -1962 -172 -1946 -155
rect -1486 -155 -1316 -138
rect -1258 -138 -458 -100
rect -1258 -155 -1088 -138
rect -1486 -172 -1470 -155
rect -1962 -188 -1470 -172
rect -1104 -172 -1088 -155
rect -628 -155 -458 -138
rect -400 -138 400 -100
rect -400 -155 -230 -138
rect -628 -172 -612 -155
rect -1104 -188 -612 -172
rect -246 -172 -230 -155
rect 230 -155 400 -138
rect 458 -138 1258 -100
rect 458 -155 628 -138
rect 230 -172 246 -155
rect -246 -188 246 -172
rect 612 -172 628 -155
rect 1088 -155 1258 -138
rect 1316 -138 2116 -100
rect 1316 -155 1486 -138
rect 1088 -172 1104 -155
rect 612 -188 1104 -172
rect 1470 -172 1486 -155
rect 1946 -155 2116 -138
rect 2174 -138 2974 -100
rect 2174 -155 2344 -138
rect 1946 -172 1962 -155
rect 1470 -188 1962 -172
rect 2328 -172 2344 -155
rect 2804 -155 2974 -138
rect 3032 -138 3832 -100
rect 3032 -155 3202 -138
rect 2804 -172 2820 -155
rect 2328 -188 2820 -172
rect 3186 -172 3202 -155
rect 3662 -155 3832 -138
rect 3662 -172 3678 -155
rect 3186 -188 3678 -172
<< polycont >>
rect -3662 138 -3202 172
rect -2804 138 -2344 172
rect -1946 138 -1486 172
rect -1088 138 -628 172
rect -230 138 230 172
rect 628 138 1088 172
rect 1486 138 1946 172
rect 2344 138 2804 172
rect 3202 138 3662 172
rect -3662 -172 -3202 -138
rect -2804 -172 -2344 -138
rect -1946 -172 -1486 -138
rect -1088 -172 -628 -138
rect -230 -172 230 -138
rect 628 -172 1088 -138
rect 1486 -172 1946 -138
rect 2344 -172 2804 -138
rect 3202 -172 3662 -138
<< locali >>
rect -3678 138 -3662 172
rect -3202 138 -3186 172
rect -2820 138 -2804 172
rect -2344 138 -2328 172
rect -1962 138 -1946 172
rect -1486 138 -1470 172
rect -1104 138 -1088 172
rect -628 138 -612 172
rect -246 138 -230 172
rect 230 138 246 172
rect 612 138 628 172
rect 1088 138 1104 172
rect 1470 138 1486 172
rect 1946 138 1962 172
rect 2328 138 2344 172
rect 2804 138 2820 172
rect 3186 138 3202 172
rect 3662 138 3678 172
rect -3878 88 -3844 104
rect -3878 -104 -3844 -88
rect -3020 88 -2986 104
rect -3020 -104 -2986 -88
rect -2162 88 -2128 104
rect -2162 -104 -2128 -88
rect -1304 88 -1270 104
rect -1304 -104 -1270 -88
rect -446 88 -412 104
rect -446 -104 -412 -88
rect 412 88 446 104
rect 412 -104 446 -88
rect 1270 88 1304 104
rect 1270 -104 1304 -88
rect 2128 88 2162 104
rect 2128 -104 2162 -88
rect 2986 88 3020 104
rect 2986 -104 3020 -88
rect 3844 88 3878 104
rect 3844 -104 3878 -88
rect -3678 -172 -3662 -138
rect -3202 -172 -3186 -138
rect -2820 -172 -2804 -138
rect -2344 -172 -2328 -138
rect -1962 -172 -1946 -138
rect -1486 -172 -1470 -138
rect -1104 -172 -1088 -138
rect -628 -172 -612 -138
rect -246 -172 -230 -138
rect 230 -172 246 -138
rect 612 -172 628 -138
rect 1088 -172 1104 -138
rect 1470 -172 1486 -138
rect 1946 -172 1962 -138
rect 2328 -172 2344 -138
rect 2804 -172 2820 -138
rect 3186 -172 3202 -138
rect 3662 -172 3678 -138
<< viali >>
rect -3624 138 -3240 172
rect -2766 138 -2382 172
rect -1908 138 -1524 172
rect -1050 138 -666 172
rect -192 138 192 172
rect 666 138 1050 172
rect 1524 138 1908 172
rect 2382 138 2766 172
rect 3240 138 3624 172
rect -3878 -88 -3844 88
rect -3020 -88 -2986 88
rect -2162 -88 -2128 88
rect -1304 -88 -1270 88
rect -446 -88 -412 88
rect 412 -88 446 88
rect 1270 -88 1304 88
rect 2128 -88 2162 88
rect 2986 -88 3020 88
rect 3844 -88 3878 88
rect -3624 -172 -3240 -138
rect -2766 -172 -2382 -138
rect -1908 -172 -1524 -138
rect -1050 -172 -666 -138
rect -192 -172 192 -138
rect 666 -172 1050 -138
rect 1524 -172 1908 -138
rect 2382 -172 2766 -138
rect 3240 -172 3624 -138
<< metal1 >>
rect -3636 172 -3228 178
rect -3636 138 -3624 172
rect -3240 138 -3228 172
rect -3636 132 -3228 138
rect -2778 172 -2370 178
rect -2778 138 -2766 172
rect -2382 138 -2370 172
rect -2778 132 -2370 138
rect -1920 172 -1512 178
rect -1920 138 -1908 172
rect -1524 138 -1512 172
rect -1920 132 -1512 138
rect -1062 172 -654 178
rect -1062 138 -1050 172
rect -666 138 -654 172
rect -1062 132 -654 138
rect -204 172 204 178
rect -204 138 -192 172
rect 192 138 204 172
rect -204 132 204 138
rect 654 172 1062 178
rect 654 138 666 172
rect 1050 138 1062 172
rect 654 132 1062 138
rect 1512 172 1920 178
rect 1512 138 1524 172
rect 1908 138 1920 172
rect 1512 132 1920 138
rect 2370 172 2778 178
rect 2370 138 2382 172
rect 2766 138 2778 172
rect 2370 132 2778 138
rect 3228 172 3636 178
rect 3228 138 3240 172
rect 3624 138 3636 172
rect 3228 132 3636 138
rect -3884 88 -3838 100
rect -3884 -88 -3878 88
rect -3844 -88 -3838 88
rect -3884 -100 -3838 -88
rect -3026 88 -2980 100
rect -3026 -88 -3020 88
rect -2986 -88 -2980 88
rect -3026 -100 -2980 -88
rect -2168 88 -2122 100
rect -2168 -88 -2162 88
rect -2128 -88 -2122 88
rect -2168 -100 -2122 -88
rect -1310 88 -1264 100
rect -1310 -88 -1304 88
rect -1270 -88 -1264 88
rect -1310 -100 -1264 -88
rect -452 88 -406 100
rect -452 -88 -446 88
rect -412 -88 -406 88
rect -452 -100 -406 -88
rect 406 88 452 100
rect 406 -88 412 88
rect 446 -88 452 88
rect 406 -100 452 -88
rect 1264 88 1310 100
rect 1264 -88 1270 88
rect 1304 -88 1310 88
rect 1264 -100 1310 -88
rect 2122 88 2168 100
rect 2122 -88 2128 88
rect 2162 -88 2168 88
rect 2122 -100 2168 -88
rect 2980 88 3026 100
rect 2980 -88 2986 88
rect 3020 -88 3026 88
rect 2980 -100 3026 -88
rect 3838 88 3884 100
rect 3838 -88 3844 88
rect 3878 -88 3884 88
rect 3838 -100 3884 -88
rect -3636 -138 -3228 -132
rect -3636 -172 -3624 -138
rect -3240 -172 -3228 -138
rect -3636 -178 -3228 -172
rect -2778 -138 -2370 -132
rect -2778 -172 -2766 -138
rect -2382 -172 -2370 -138
rect -2778 -178 -2370 -172
rect -1920 -138 -1512 -132
rect -1920 -172 -1908 -138
rect -1524 -172 -1512 -138
rect -1920 -178 -1512 -172
rect -1062 -138 -654 -132
rect -1062 -172 -1050 -138
rect -666 -172 -654 -138
rect -1062 -178 -654 -172
rect -204 -138 204 -132
rect -204 -172 -192 -138
rect 192 -172 204 -138
rect -204 -178 204 -172
rect 654 -138 1062 -132
rect 654 -172 666 -138
rect 1050 -172 1062 -138
rect 654 -178 1062 -172
rect 1512 -138 1920 -132
rect 1512 -172 1524 -138
rect 1908 -172 1920 -138
rect 1512 -178 1920 -172
rect 2370 -138 2778 -132
rect 2370 -172 2382 -138
rect 2766 -172 2778 -138
rect 2370 -178 2778 -172
rect 3228 -138 3636 -132
rect 3228 -172 3240 -138
rect 3624 -172 3636 -138
rect 3228 -178 3636 -172
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 1 l 4 m 1 nf 9 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>

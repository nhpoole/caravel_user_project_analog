magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nmos >>
rect -745 -200 -545 200
rect -487 -200 -287 200
rect -229 -200 -29 200
rect 29 -200 229 200
rect 287 -200 487 200
rect 545 -200 745 200
<< ndiff >>
rect -803 188 -745 200
rect -803 -188 -791 188
rect -757 -188 -745 188
rect -803 -200 -745 -188
rect -545 188 -487 200
rect -545 -188 -533 188
rect -499 -188 -487 188
rect -545 -200 -487 -188
rect -287 188 -229 200
rect -287 -188 -275 188
rect -241 -188 -229 188
rect -287 -200 -229 -188
rect -29 188 29 200
rect -29 -188 -17 188
rect 17 -188 29 188
rect -29 -200 29 -188
rect 229 188 287 200
rect 229 -188 241 188
rect 275 -188 287 188
rect 229 -200 287 -188
rect 487 188 545 200
rect 487 -188 499 188
rect 533 -188 545 188
rect 487 -200 545 -188
rect 745 188 803 200
rect 745 -188 757 188
rect 791 -188 803 188
rect 745 -200 803 -188
<< ndiffc >>
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
<< poly >>
rect -711 272 -579 288
rect -711 255 -695 272
rect -745 238 -695 255
rect -595 255 -579 272
rect -453 272 -321 288
rect -453 255 -437 272
rect -595 238 -545 255
rect -745 200 -545 238
rect -487 238 -437 255
rect -337 255 -321 272
rect -195 272 -63 288
rect -195 255 -179 272
rect -337 238 -287 255
rect -487 200 -287 238
rect -229 238 -179 255
rect -79 255 -63 272
rect 63 272 195 288
rect 63 255 79 272
rect -79 238 -29 255
rect -229 200 -29 238
rect 29 238 79 255
rect 179 255 195 272
rect 321 272 453 288
rect 321 255 337 272
rect 179 238 229 255
rect 29 200 229 238
rect 287 238 337 255
rect 437 255 453 272
rect 579 272 711 288
rect 579 255 595 272
rect 437 238 487 255
rect 287 200 487 238
rect 545 238 595 255
rect 695 255 711 272
rect 695 238 745 255
rect 545 200 745 238
rect -745 -238 -545 -200
rect -745 -255 -695 -238
rect -711 -272 -695 -255
rect -595 -255 -545 -238
rect -487 -238 -287 -200
rect -487 -255 -437 -238
rect -595 -272 -579 -255
rect -711 -288 -579 -272
rect -453 -272 -437 -255
rect -337 -255 -287 -238
rect -229 -238 -29 -200
rect -229 -255 -179 -238
rect -337 -272 -321 -255
rect -453 -288 -321 -272
rect -195 -272 -179 -255
rect -79 -255 -29 -238
rect 29 -238 229 -200
rect 29 -255 79 -238
rect -79 -272 -63 -255
rect -195 -288 -63 -272
rect 63 -272 79 -255
rect 179 -255 229 -238
rect 287 -238 487 -200
rect 287 -255 337 -238
rect 179 -272 195 -255
rect 63 -288 195 -272
rect 321 -272 337 -255
rect 437 -255 487 -238
rect 545 -238 745 -200
rect 545 -255 595 -238
rect 437 -272 453 -255
rect 321 -288 453 -272
rect 579 -272 595 -255
rect 695 -255 745 -238
rect 695 -272 711 -255
rect 579 -288 711 -272
<< polycont >>
rect -695 238 -595 272
rect -437 238 -337 272
rect -179 238 -79 272
rect 79 238 179 272
rect 337 238 437 272
rect 595 238 695 272
rect -695 -272 -595 -238
rect -437 -272 -337 -238
rect -179 -272 -79 -238
rect 79 -272 179 -238
rect 337 -272 437 -238
rect 595 -272 695 -238
<< locali >>
rect -711 238 -695 272
rect -595 238 -579 272
rect -453 238 -437 272
rect -337 238 -321 272
rect -195 238 -179 272
rect -79 238 -63 272
rect 63 238 79 272
rect 179 238 195 272
rect 321 238 337 272
rect 437 238 453 272
rect 579 238 595 272
rect 695 238 711 272
rect -791 188 -757 204
rect -791 -204 -757 -188
rect -533 188 -499 204
rect -533 -204 -499 -188
rect -275 188 -241 204
rect -275 -204 -241 -188
rect -17 188 17 204
rect -17 -204 17 -188
rect 241 188 275 204
rect 241 -204 275 -188
rect 499 188 533 204
rect 499 -204 533 -188
rect 757 188 791 204
rect 757 -204 791 -188
rect -711 -272 -695 -238
rect -595 -272 -579 -238
rect -453 -272 -437 -238
rect -337 -272 -321 -238
rect -195 -272 -179 -238
rect -79 -272 -63 -238
rect 63 -272 79 -238
rect 179 -272 195 -238
rect 321 -272 337 -238
rect 437 -272 453 -238
rect 579 -272 595 -238
rect 695 -272 711 -238
<< viali >>
rect -687 238 -603 272
rect -429 238 -345 272
rect -171 238 -87 272
rect 87 238 171 272
rect 345 238 429 272
rect 603 238 687 272
rect -791 -188 -757 188
rect -533 -188 -499 188
rect -275 -188 -241 188
rect -17 -188 17 188
rect 241 -188 275 188
rect 499 -188 533 188
rect 757 -188 791 188
rect -687 -272 -603 -238
rect -429 -272 -345 -238
rect -171 -272 -87 -238
rect 87 -272 171 -238
rect 345 -272 429 -238
rect 603 -272 687 -238
<< metal1 >>
rect -699 272 -591 278
rect -699 238 -687 272
rect -603 238 -591 272
rect -699 232 -591 238
rect -441 272 -333 278
rect -441 238 -429 272
rect -345 238 -333 272
rect -441 232 -333 238
rect -183 272 -75 278
rect -183 238 -171 272
rect -87 238 -75 272
rect -183 232 -75 238
rect 75 272 183 278
rect 75 238 87 272
rect 171 238 183 272
rect 75 232 183 238
rect 333 272 441 278
rect 333 238 345 272
rect 429 238 441 272
rect 333 232 441 238
rect 591 272 699 278
rect 591 238 603 272
rect 687 238 699 272
rect 591 232 699 238
rect -797 188 -751 200
rect -797 -188 -791 188
rect -757 -188 -751 188
rect -797 -200 -751 -188
rect -539 188 -493 200
rect -539 -188 -533 188
rect -499 -188 -493 188
rect -539 -200 -493 -188
rect -281 188 -235 200
rect -281 -188 -275 188
rect -241 -188 -235 188
rect -281 -200 -235 -188
rect -23 188 23 200
rect -23 -188 -17 188
rect 17 -188 23 188
rect -23 -200 23 -188
rect 235 188 281 200
rect 235 -188 241 188
rect 275 -188 281 188
rect 235 -200 281 -188
rect 493 188 539 200
rect 493 -188 499 188
rect 533 -188 539 188
rect 493 -200 539 -188
rect 751 188 797 200
rect 751 -188 757 188
rect 791 -188 797 188
rect 751 -200 797 -188
rect -699 -238 -591 -232
rect -699 -272 -687 -238
rect -603 -272 -591 -238
rect -699 -278 -591 -272
rect -441 -238 -333 -232
rect -441 -272 -429 -238
rect -345 -272 -333 -238
rect -441 -278 -333 -272
rect -183 -238 -75 -232
rect -183 -272 -171 -238
rect -87 -272 -75 -238
rect -183 -278 -75 -272
rect 75 -238 183 -232
rect 75 -272 87 -238
rect 171 -272 183 -238
rect 75 -278 183 -272
rect 333 -238 441 -232
rect 333 -272 345 -238
rect 429 -272 441 -238
rect 333 -278 441 -272
rect 591 -238 699 -232
rect 591 -272 603 -238
rect 687 -272 699 -238
rect 591 -278 699 -272
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string parameters w 2 l 1 m 1 nf 6 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< metal3 >>
rect -1150 -1100 1050 1100
<< mimcap >>
rect -1050 960 950 1000
rect -1050 -960 -1010 960
rect 910 -960 950 960
rect -1050 -1000 950 -960
<< mimcapcontact >>
rect -1010 -960 910 960
<< metal4 >>
rect -1011 960 911 961
rect -1011 -960 -1010 960
rect 910 -960 911 960
rect -1011 -961 911 -960
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -1150 -1100 1050 1100
string parameters w 10.00 l 10.00 val 207.6 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
string library sky130
<< end >>

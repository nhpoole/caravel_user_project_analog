magic
tech sky130A
magscale 1 2
timestamp 1624302123
<< nwell >>
rect 97364 586526 98856 587312
<< metal1 >>
rect 171904 702110 172024 702118
rect 171904 701994 171906 702110
rect 172022 701994 172024 702110
rect 171904 701868 172024 701994
rect 174410 702110 174530 702118
rect 174410 701994 174412 702110
rect 174528 701994 174530 702110
rect 174410 701868 174530 701994
rect 223692 702110 223812 702118
rect 223692 701994 223694 702110
rect 223810 701994 223812 702110
rect 223692 701868 223812 701994
rect 226092 702110 226212 702118
rect 226092 701994 226094 702110
rect 226210 701994 226212 702110
rect 226092 701868 226212 701994
rect 325330 702110 325450 702118
rect 325330 701994 325332 702110
rect 325448 701994 325450 702110
rect 325330 701868 325450 701994
rect 327840 702110 327960 702118
rect 327840 701994 327842 702110
rect 327958 701994 327960 702110
rect 327840 701868 327960 701994
rect 171904 701148 172024 701262
rect 171904 701032 171906 701148
rect 172022 701032 172024 701148
rect 171904 701024 172024 701032
rect 174410 701148 174530 701262
rect 174410 701032 174412 701148
rect 174528 701032 174530 701148
rect 174410 701024 174530 701032
rect 223692 701148 223812 701262
rect 223692 701032 223694 701148
rect 223810 701032 223812 701148
rect 223692 701024 223812 701032
rect 226092 701148 226212 701262
rect 226092 701032 226094 701148
rect 226210 701032 226212 701148
rect 226092 701024 226212 701032
rect 325330 701148 325450 701262
rect 325330 701032 325332 701148
rect 325448 701032 325450 701148
rect 325330 701024 325450 701032
rect 327840 701148 327960 701262
rect 327840 701032 327842 701148
rect 327958 701032 327960 701148
rect 327840 701024 327960 701032
rect 281522 638598 281582 638604
rect 281050 638594 281582 638598
rect 281050 638542 281526 638594
rect 281578 638542 281582 638594
rect 281050 638538 281582 638542
rect 281522 638532 281582 638538
rect 270574 595388 270674 595394
rect 271642 595388 271742 595394
rect 270574 595364 271742 595388
rect 270574 595312 270598 595364
rect 270650 595312 271666 595364
rect 271718 595312 271742 595364
rect 270574 595288 271742 595312
rect 270574 595282 270674 595288
rect 271642 595282 271742 595288
rect 251483 554476 251773 554522
rect 579046 14659 579299 14662
rect 579046 14543 579055 14659
rect 579171 14543 579299 14659
rect 579046 14542 579299 14543
rect 579899 14659 580271 14662
rect 579899 14543 580146 14659
rect 580262 14543 580271 14659
rect 579899 14542 580271 14543
rect 579046 14540 579267 14542
rect 579928 14540 580271 14542
rect 579058 9933 579311 9936
rect 579058 9817 579067 9933
rect 579183 9817 579311 9933
rect 579058 9816 579311 9817
rect 579911 9933 580283 9936
rect 579911 9817 580158 9933
rect 580274 9817 580283 9933
rect 579911 9816 580283 9817
rect 579058 9814 579279 9816
rect 579940 9814 580283 9816
rect 579170 5203 579391 5206
rect 579170 5087 579179 5203
rect 579295 5087 579391 5203
rect 579170 5084 579391 5087
rect 580052 5203 580395 5206
rect 580052 5087 580270 5203
rect 580386 5087 580395 5203
rect 580052 5084 580395 5087
<< via1 >>
rect 171906 701994 172022 702110
rect 174412 701994 174528 702110
rect 223694 701994 223810 702110
rect 226094 701994 226210 702110
rect 325332 701994 325448 702110
rect 327842 701994 327958 702110
rect 171906 701032 172022 701148
rect 174412 701032 174528 701148
rect 223694 701032 223810 701148
rect 226094 701032 226210 701148
rect 325332 701032 325448 701148
rect 327842 701032 327958 701148
rect 281526 638542 281578 638594
rect 270598 595312 270650 595364
rect 271666 595312 271718 595364
rect 579055 14543 579171 14659
rect 580146 14543 580262 14659
rect 579067 9817 579183 9933
rect 580158 9817 580274 9933
rect 579179 5087 579295 5203
rect 580270 5087 580386 5203
<< metal2 >>
rect 171904 702112 172024 702121
rect 174410 702112 174530 702121
rect 223692 702112 223812 702121
rect 226092 702112 226212 702121
rect 325330 702112 325450 702121
rect 327840 702112 327960 702121
rect 171898 702110 172030 702112
rect 171898 701994 171906 702110
rect 172022 701994 172030 702110
rect 171898 701992 172030 701994
rect 174404 702110 174536 702112
rect 174404 701994 174412 702110
rect 174528 701994 174536 702110
rect 174404 701992 174536 701994
rect 223686 702110 223818 702112
rect 223686 701994 223694 702110
rect 223810 701994 223818 702110
rect 223686 701992 223818 701994
rect 226086 702110 226218 702112
rect 226086 701994 226094 702110
rect 226210 701994 226218 702110
rect 226086 701992 226218 701994
rect 325324 702110 325456 702112
rect 325324 701994 325332 702110
rect 325448 701994 325456 702110
rect 325324 701992 325456 701994
rect 327834 702110 327966 702112
rect 327834 701994 327842 702110
rect 327958 701994 327966 702110
rect 327834 701992 327966 701994
rect 171904 701983 172024 701992
rect 174410 701983 174530 701992
rect 223692 701983 223812 701992
rect 226092 701983 226212 701992
rect 325330 701983 325450 701992
rect 327840 701983 327960 701992
rect 128656 701378 134915 701804
rect 26120 700682 26580 700691
rect 24004 700680 26580 700682
rect 24004 700224 26122 700680
rect 26578 700224 26580 700680
rect 24004 700222 26580 700224
rect 26120 700213 26580 700222
rect 69181 700256 73612 700674
rect 18310 697685 18730 697689
rect 18305 697658 20597 697685
rect 18305 697282 18332 697658
rect 18708 697282 20597 697658
rect 28697 697645 29117 697649
rect 18305 697255 20597 697282
rect 24191 697618 29122 697645
rect 18310 697251 18730 697255
rect 24191 697242 28719 697618
rect 29095 697242 29122 697618
rect 24191 697215 29122 697242
rect 28697 697211 29117 697215
rect 12317 694671 30612 694688
rect 12317 694295 30210 694671
rect 30586 694295 30612 694671
rect 12317 694278 30612 694295
rect 7656 685938 10141 685950
rect 7656 685562 9744 685938
rect 10120 685562 10141 685938
rect 7656 685550 10141 685562
rect 10111 683066 11033 683071
rect 2919 682855 3223 682859
rect 2914 682846 4271 682855
rect 2914 682550 2923 682846
rect 3219 682550 4271 682846
rect 2914 682541 4271 682550
rect 2919 682537 3223 682541
rect 7828 682498 11033 683066
rect 9010 679962 9410 679975
rect 7544 679954 9410 679962
rect 7544 679578 9022 679954
rect 9398 679578 9410 679954
rect 7544 679570 9410 679578
rect 9010 679557 9410 679570
rect 10111 678139 11033 682498
rect 12317 679971 12727 694278
rect 69181 690560 69599 700256
rect 133170 699222 133538 699267
rect 133170 698926 133206 699222
rect 133502 698926 133538 699222
rect 130731 698878 131181 698882
rect 122377 698862 122827 698866
rect 122372 698820 125904 698862
rect 122372 698444 122414 698820
rect 122790 698444 125904 698820
rect 122372 698402 125904 698444
rect 129100 698836 131186 698878
rect 129100 698460 130768 698836
rect 131144 698460 131186 698836
rect 129100 698418 131186 698460
rect 130731 698414 131181 698418
rect 122377 698398 122827 698402
rect 70569 697684 70947 697688
rect 70564 697678 73834 697684
rect 70564 697302 70570 697678
rect 70946 697302 73834 697678
rect 70564 697296 73834 697302
rect 77192 697662 79362 697668
rect 77192 697652 79367 697662
rect 70569 697292 70947 697296
rect 77192 697280 78990 697652
rect 78989 697276 78990 697280
rect 79366 697276 79367 697652
rect 78989 697266 79367 697276
rect 81976 695830 82400 695845
rect 81976 695454 82000 695830
rect 82376 695454 82400 695830
rect 133170 695774 133538 698926
rect 81976 695439 82400 695454
rect 122457 695738 133538 695774
rect 122457 695442 122502 695738
rect 122798 695442 133538 695738
rect 81985 694670 82391 695439
rect 122457 695406 133538 695442
rect 71588 694655 82391 694670
rect 71588 694279 71612 694655
rect 71988 694279 82391 694655
rect 71588 694264 82391 694279
rect 69181 690184 69202 690560
rect 69578 690184 69599 690560
rect 69181 690154 69599 690184
rect 134489 690566 134915 701378
rect 171898 701148 172030 701150
rect 171898 701032 171906 701148
rect 172022 701032 172030 701148
rect 171898 701030 172030 701032
rect 174404 701148 174536 701150
rect 174404 701032 174412 701148
rect 174528 701032 174536 701148
rect 174404 701030 174536 701032
rect 223686 701148 223818 701150
rect 223686 701032 223694 701148
rect 223810 701032 223818 701148
rect 223686 701030 223818 701032
rect 226086 701148 226218 701150
rect 226086 701032 226094 701148
rect 226210 701032 226218 701148
rect 226086 701030 226218 701032
rect 325324 701148 325456 701150
rect 325324 701032 325332 701148
rect 325448 701032 325456 701148
rect 325324 701030 325456 701032
rect 327834 701148 327966 701150
rect 327834 701032 327842 701148
rect 327958 701032 327966 701148
rect 327834 701030 327966 701032
rect 171904 699140 172024 701030
rect 174410 700926 174530 701030
rect 223692 700926 223812 701030
rect 226092 700926 226212 701030
rect 325330 700926 325450 701030
rect 171895 699108 172033 699140
rect 171895 699052 171936 699108
rect 171992 699052 172033 699108
rect 171895 699020 172033 699052
rect 174410 699110 174514 700926
rect 196531 700814 197131 700837
rect 196531 700278 196563 700814
rect 197099 700278 197131 700814
rect 219622 700323 220106 700328
rect 196531 700255 197131 700278
rect 219618 700314 220110 700323
rect 174410 699054 174434 699110
rect 174490 699054 174514 699110
rect 174410 699021 174514 699054
rect 194103 697888 194581 697890
rect 194103 697432 194114 697888
rect 194570 697432 194581 697888
rect 194103 697430 194581 697432
rect 186408 695448 186788 695500
rect 186399 695446 186797 695448
rect 186399 695070 186410 695446
rect 186786 695070 186797 695446
rect 186399 695068 186797 695070
rect 185235 694628 185397 694632
rect 185235 694492 185248 694628
rect 185384 694492 185397 694628
rect 185235 694488 185397 694492
rect 134489 690190 134514 690566
rect 134890 690190 134915 690566
rect 134489 690156 134915 690190
rect 12308 679954 12736 679971
rect 12308 679578 12334 679954
rect 12710 679578 12736 679954
rect 12308 679561 12736 679578
rect 7576 677217 11033 678139
rect 4122 657477 5114 657482
rect 4118 657454 5118 657477
rect 4118 656518 4150 657454
rect 5086 656518 5118 657454
rect 4118 656495 5118 656518
rect 4122 338726 5114 656495
rect 7576 549431 8498 677217
rect 9587 659438 10507 659461
rect 9587 658582 9619 659438
rect 10475 658582 10507 659438
rect 9587 658559 10507 658582
rect 7576 549135 7870 549431
rect 8166 549135 8498 549431
rect 7576 549052 8498 549135
rect 9596 600628 10498 658559
rect 11758 655201 12658 655206
rect 11754 655184 12662 655201
rect 11754 654328 11780 655184
rect 12636 654328 12662 655184
rect 11754 654311 12662 654328
rect 9596 600492 9926 600628
rect 10062 600492 10498 600628
rect 4122 338670 4626 338726
rect 4682 338670 5114 338726
rect 4122 338630 5114 338670
rect 6634 548692 7768 548794
rect 6634 548396 7102 548692
rect 7398 548396 7768 548692
rect 6634 81638 7768 548396
rect 9596 547542 10498 600492
rect 9596 547326 9980 547542
rect 10196 547326 10498 547542
rect 9596 121314 10498 547326
rect 11758 381948 12658 654311
rect 91824 638532 94332 638644
rect 90749 622150 90827 622152
rect 90749 622136 90760 622150
rect 90570 622108 90760 622136
rect 90749 622094 90760 622108
rect 90816 622094 90827 622150
rect 90749 622092 90827 622094
rect 90665 619974 90743 619976
rect 90665 619960 90676 619974
rect 90574 619932 90676 619960
rect 90665 619918 90676 619932
rect 90732 619918 90743 619974
rect 90665 619916 90743 619918
rect 90953 617730 91031 617732
rect 90953 617716 90964 617730
rect 90574 617688 90964 617716
rect 90953 617674 90964 617688
rect 91020 617674 91031 617730
rect 90953 617672 91031 617674
rect 90751 615486 90829 615488
rect 90751 615472 90762 615486
rect 90570 615444 90762 615472
rect 90751 615430 90762 615444
rect 90818 615430 90829 615486
rect 90751 615428 90829 615430
rect 90741 613242 90819 613244
rect 90741 613228 90752 613242
rect 90574 613200 90752 613228
rect 90741 613186 90752 613200
rect 90808 613186 90819 613242
rect 90741 613184 90819 613186
rect 90699 611066 90777 611068
rect 90699 611052 90710 611066
rect 90572 611024 90710 611052
rect 90699 611010 90710 611024
rect 90766 611010 90777 611066
rect 90699 611008 90777 611010
rect 90723 608822 90801 608824
rect 90723 608808 90734 608822
rect 90574 608780 90734 608808
rect 90723 608766 90734 608780
rect 90790 608766 90801 608822
rect 90723 608764 90801 608766
rect 90657 606578 90735 606580
rect 90657 606564 90668 606578
rect 90572 606536 90668 606564
rect 90657 606522 90668 606536
rect 90724 606522 90735 606578
rect 90657 606520 90735 606522
rect 90691 604334 90769 604336
rect 90691 604320 90702 604334
rect 90570 604292 90702 604320
rect 90691 604278 90702 604292
rect 90758 604278 90769 604334
rect 90691 604276 90769 604278
rect 74050 602048 74542 602076
rect 11758 381892 12260 381948
rect 12316 381892 12658 381948
rect 11758 381792 12658 381892
rect 14310 601324 14978 601382
rect 14310 601188 14610 601324
rect 14746 601188 14978 601324
rect 14310 550244 14978 601188
rect 14310 550028 14590 550244
rect 14806 550028 14978 550244
rect 14310 248936 14978 550028
rect 16692 596943 17468 596986
rect 16692 596647 16920 596943
rect 17216 596647 17468 596943
rect 16692 468392 17468 596647
rect 74050 594530 74167 602048
rect 74718 601282 74746 602076
rect 74693 601280 74771 601282
rect 74693 601224 74704 601280
rect 74760 601224 74771 601280
rect 74693 601222 74771 601224
rect 82538 600586 82566 602082
rect 90358 601720 90386 602162
rect 91824 602118 91936 638532
rect 98678 619968 98798 620009
rect 98678 619912 98710 619968
rect 98766 619912 98798 619968
rect 98365 617746 98483 617786
rect 98365 617690 98396 617746
rect 98452 617690 98483 617746
rect 98061 615490 98179 615530
rect 98061 615434 98092 615490
rect 98148 615434 98179 615490
rect 97757 613232 97875 613272
rect 97757 613176 97788 613232
rect 97844 613176 97875 613232
rect 97467 611024 97585 611064
rect 97467 610968 97498 611024
rect 97554 610968 97585 611024
rect 97187 608826 97305 608866
rect 97187 608770 97218 608826
rect 97274 608770 97305 608826
rect 96883 606570 97001 606610
rect 96883 606514 96914 606570
rect 96970 606514 97001 606570
rect 90738 602076 91936 602118
rect 90570 602048 91936 602076
rect 90738 602006 91936 602048
rect 82513 600584 82591 600586
rect 82513 600528 82524 600584
rect 82580 600528 82591 600584
rect 82513 600526 82591 600528
rect 74050 594474 74080 594530
rect 74136 594474 74167 594530
rect 74050 594435 74167 594474
rect 90315 578416 90430 601720
rect 91824 596824 91936 602006
rect 91824 596768 91852 596824
rect 91908 596768 91936 596824
rect 91824 596731 91936 596768
rect 96629 604336 96747 604376
rect 96629 604280 96660 604336
rect 96716 604280 96747 604336
rect 96629 594258 96747 604280
rect 96625 594232 96751 594258
rect 96625 594176 96660 594232
rect 96716 594176 96751 594232
rect 96625 594150 96751 594176
rect 96629 594145 96747 594150
rect 96883 593962 97001 606514
rect 96879 593936 97005 593962
rect 96879 593880 96914 593936
rect 96970 593880 97005 593936
rect 96879 593854 97005 593880
rect 96883 593849 97001 593854
rect 97187 593694 97305 608770
rect 97183 593668 97309 593694
rect 97183 593612 97218 593668
rect 97274 593612 97309 593668
rect 97183 593586 97309 593612
rect 97187 593581 97305 593586
rect 97467 593424 97585 610968
rect 97463 593398 97589 593424
rect 97463 593342 97498 593398
rect 97554 593342 97589 593398
rect 97463 593316 97589 593342
rect 97467 593311 97585 593316
rect 97757 593112 97875 613176
rect 97753 593086 97879 593112
rect 97753 593030 97788 593086
rect 97844 593030 97879 593086
rect 97753 593004 97879 593030
rect 97757 592999 97875 593004
rect 98061 592822 98179 615434
rect 98057 592796 98183 592822
rect 98057 592740 98092 592796
rect 98148 592740 98183 592796
rect 98057 592714 98183 592740
rect 98061 592709 98179 592714
rect 98365 592532 98483 617690
rect 98361 592506 98487 592532
rect 98361 592450 98396 592506
rect 98452 592450 98487 592506
rect 98361 592424 98487 592450
rect 98365 592419 98483 592424
rect 98678 592263 98798 619912
rect 185244 617670 185388 694488
rect 185649 693166 185658 693302
rect 185794 693166 185803 693302
rect 185244 617614 185288 617670
rect 185344 617614 185388 617670
rect 185244 617570 185388 617614
rect 185658 617656 185794 693166
rect 186408 617739 186788 695068
rect 194112 633070 194572 697430
rect 196540 689907 197122 700255
rect 219618 699858 219636 700314
rect 220092 699858 220110 700314
rect 219618 699849 220110 699858
rect 209714 698010 213770 698398
rect 209714 693983 210102 698010
rect 219622 695486 220106 699849
rect 210649 695448 211019 695452
rect 210644 695406 213252 695448
rect 210644 695110 210686 695406
rect 210982 695110 213252 695406
rect 210644 695068 213252 695110
rect 210649 695064 211019 695068
rect 217014 695002 220106 695486
rect 221404 699222 221768 699265
rect 221404 698926 221438 699222
rect 221734 698926 221768 699222
rect 223696 699124 223800 700926
rect 223696 699068 223720 699124
rect 223776 699068 223800 699124
rect 223696 699035 223800 699068
rect 226094 699144 226198 700926
rect 321254 700815 321929 700820
rect 313064 700809 313742 700814
rect 313060 700783 313746 700809
rect 264679 700460 264881 700484
rect 264679 700324 264712 700460
rect 264848 700324 264881 700460
rect 264679 700300 264881 700324
rect 226094 699088 226118 699144
rect 226174 699088 226198 699144
rect 226094 699055 226198 699088
rect 202378 693968 210102 693983
rect 202378 693593 209720 693968
rect 202378 692802 202768 693593
rect 209714 693592 209720 693593
rect 210096 693592 210102 693968
rect 209714 693577 210102 693592
rect 201658 692412 202768 692802
rect 204962 692393 205298 692397
rect 204957 692368 214309 692393
rect 221404 692392 221768 698926
rect 204957 692072 204982 692368
rect 205278 692072 214309 692368
rect 204957 692047 214309 692072
rect 204962 692043 205298 692047
rect 216576 692028 221768 692392
rect 196540 689325 198199 689907
rect 201703 689341 203819 689923
rect 201328 686779 202816 686804
rect 201328 686483 202486 686779
rect 202782 686483 202816 686779
rect 201328 686458 202816 686483
rect 203237 684908 203819 689341
rect 196540 684326 203819 684908
rect 196540 643266 197122 684326
rect 264688 659432 264872 700300
rect 313060 700167 313095 700783
rect 313711 700167 313746 700783
rect 313060 700141 313746 700167
rect 321250 700790 321933 700815
rect 321250 700174 321283 700790
rect 321899 700174 321933 700790
rect 321250 700150 321933 700174
rect 310798 699220 311178 699253
rect 310798 698924 310840 699220
rect 311136 698924 311178 699220
rect 310798 698891 311178 698924
rect 310807 692004 311169 698891
rect 313064 695177 313742 700141
rect 314732 698040 315200 698049
rect 314732 698034 316514 698040
rect 314732 697578 314738 698034
rect 315194 697578 316514 698034
rect 314732 697572 316514 697578
rect 314732 697563 315200 697572
rect 313064 694499 316479 695177
rect 321254 695160 321929 700150
rect 325346 699084 325450 700926
rect 325346 699028 325370 699084
rect 325426 699028 325450 699084
rect 325346 698995 325450 699028
rect 327840 700926 327960 701030
rect 327840 699096 327944 700926
rect 327840 699040 327864 699096
rect 327920 699040 327944 699096
rect 327840 699007 327944 699040
rect 401679 699560 406962 699946
rect 323703 697026 324535 697045
rect 323703 696250 323731 697026
rect 324507 696250 324535 697026
rect 323703 696231 324535 696250
rect 319471 694485 321929 695160
rect 310807 691642 316624 692004
rect 282148 663358 282320 663367
rect 282148 663222 282166 663358
rect 282302 663222 282320 663358
rect 282148 663213 282320 663222
rect 279750 661698 279828 661700
rect 279750 661642 279761 661698
rect 279817 661642 279828 661698
rect 279750 661640 279828 661642
rect 264688 659248 265668 659432
rect 215174 657014 215430 657025
rect 215174 656798 215194 657014
rect 215410 656798 215430 657014
rect 215174 656787 215430 656798
rect 196540 643206 199146 643266
rect 196540 643204 197122 643206
rect 215183 638231 215421 656787
rect 215877 654758 216147 654776
rect 215877 654542 215904 654758
rect 216120 654542 216147 654758
rect 215877 654524 216147 654542
rect 215886 638864 216138 654524
rect 222630 648426 222758 648435
rect 222630 648390 222870 648426
rect 222630 648334 222666 648390
rect 222722 648334 222870 648390
rect 222630 648298 222870 648334
rect 222630 648289 222758 648298
rect 265484 639622 265668 659248
rect 279759 657346 279819 661640
rect 282157 646930 282311 663213
rect 281522 646776 282311 646930
rect 265484 639438 266472 639622
rect 220299 638864 220389 638868
rect 215886 638842 220394 638864
rect 215886 638786 220316 638842
rect 220372 638786 220394 638842
rect 215886 638764 220394 638786
rect 220299 638760 220389 638764
rect 215183 637993 216470 638231
rect 216232 634334 216470 637993
rect 220155 634334 220245 634338
rect 216232 634312 220250 634334
rect 216232 634256 220172 634312
rect 220228 634256 220250 634312
rect 216232 634234 220250 634256
rect 216232 634233 216470 634234
rect 220155 634230 220245 634234
rect 194112 632610 202278 633070
rect 201818 631492 202278 632610
rect 201818 631432 203356 631492
rect 201818 631430 202278 631432
rect 266288 629562 266472 639438
rect 281522 638598 281582 646776
rect 294194 640108 294561 640110
rect 294194 640052 294494 640108
rect 294550 640052 294561 640108
rect 294194 640050 294561 640052
rect 281516 638594 281588 638598
rect 281516 638542 281526 638594
rect 281578 638542 281588 638594
rect 281516 638538 281588 638542
rect 285231 634098 285433 634103
rect 285227 634070 285437 634098
rect 285227 633934 285264 634070
rect 285400 633934 285437 634070
rect 285227 633906 285437 633934
rect 267168 632734 267388 632767
rect 267168 632598 267210 632734
rect 267346 632598 267388 632734
rect 267168 632565 267388 632598
rect 265750 629378 266472 629562
rect 244663 628666 244865 628690
rect 265750 628686 265934 629378
rect 244663 628530 244696 628666
rect 244832 628530 244865 628666
rect 244663 628506 244865 628530
rect 265741 628662 265943 628686
rect 265741 628526 265774 628662
rect 265910 628526 265943 628662
rect 244672 624544 244856 628506
rect 265741 628502 265943 628526
rect 245661 628324 245881 628357
rect 267177 628352 267379 632565
rect 285231 632479 285433 633906
rect 285222 632446 285442 632479
rect 285222 632310 285264 632446
rect 285400 632310 285442 632446
rect 285222 632277 285442 632310
rect 282607 631908 282725 631930
rect 289032 631925 289132 631930
rect 282607 631852 282638 631908
rect 282694 631852 282725 631908
rect 282607 631830 282725 631852
rect 289028 631908 289136 631925
rect 289028 631852 289054 631908
rect 289110 631852 289136 631908
rect 289028 631835 289136 631852
rect 289032 630778 289132 631835
rect 289032 630776 295028 630778
rect 289032 630678 295332 630776
rect 294048 630001 294304 630006
rect 294044 629986 294308 630001
rect 294044 629770 294068 629986
rect 294284 629770 294308 629986
rect 294044 629755 294308 629770
rect 291971 629454 292089 629476
rect 291971 629398 292002 629454
rect 292058 629398 292089 629454
rect 291971 629376 292089 629398
rect 245661 628188 245703 628324
rect 245839 628188 245881 628324
rect 245661 628155 245881 628188
rect 267173 628324 267383 628352
rect 267173 628188 267210 628324
rect 267346 628188 267383 628324
rect 267173 628160 267383 628188
rect 267177 628155 267379 628160
rect 245670 625724 245872 628155
rect 291980 626835 292080 629376
rect 291976 626818 292084 626835
rect 291976 626762 292002 626818
rect 292058 626762 292084 626818
rect 291976 626745 292084 626762
rect 291980 626740 292080 626745
rect 294048 625760 294304 629755
rect 294822 627029 295332 630678
rect 294813 627002 295341 627029
rect 294813 626546 294849 627002
rect 295305 626546 295341 627002
rect 294813 626519 295341 626546
rect 245670 625668 245732 625724
rect 245788 625668 245872 625724
rect 245670 625644 245872 625668
rect 294039 625740 294313 625760
rect 294039 625524 294068 625740
rect 294284 625524 294313 625740
rect 294039 625504 294313 625524
rect 292225 623746 292315 623750
rect 292220 623724 294425 623746
rect 292220 623668 292242 623724
rect 292298 623668 294338 623724
rect 294394 623668 294425 623724
rect 292220 623646 294425 623668
rect 292225 623642 292315 623646
rect 185658 617600 185698 617656
rect 185754 617600 185794 617656
rect 185658 617560 185794 617600
rect 186404 617702 186792 617739
rect 186404 617406 186450 617702
rect 186746 617406 186792 617702
rect 186404 617369 186792 617406
rect 186408 617364 186788 617369
rect 182719 615892 182837 615914
rect 182719 615836 182750 615892
rect 182806 615836 182837 615892
rect 182719 615814 182837 615836
rect 182728 605699 182828 615814
rect 183057 615486 183175 615508
rect 183057 615430 183088 615486
rect 183144 615430 183175 615486
rect 183057 615408 183175 615430
rect 183066 607683 183166 615408
rect 183062 607666 183170 607683
rect 183062 607610 183088 607666
rect 183144 607610 183170 607666
rect 183062 607593 183170 607610
rect 183066 607588 183166 607593
rect 182724 605682 182832 605699
rect 182724 605626 182750 605682
rect 182806 605626 182832 605682
rect 182724 605609 182832 605626
rect 182728 605604 182828 605609
rect 270579 595388 270669 595392
rect 271642 595388 271742 602430
rect 270568 595366 270680 595388
rect 270568 595310 270596 595366
rect 270652 595310 270680 595366
rect 270568 595288 270680 595310
rect 271636 595364 271748 595388
rect 271636 595312 271666 595364
rect 271718 595312 271748 595364
rect 271636 595288 271748 595312
rect 270579 595284 270669 595288
rect 98674 592236 98802 592263
rect 98674 592180 98710 592236
rect 98766 592180 98802 592236
rect 98674 592153 98802 592180
rect 98678 592148 98798 592153
rect 91840 587526 94346 587638
rect 90313 578391 90436 578416
rect 90313 578335 90346 578391
rect 90402 578335 90436 578391
rect 90313 578311 90436 578335
rect 90315 578299 90430 578311
rect 90681 568624 90759 568626
rect 90681 568610 90692 568624
rect 90590 568582 90692 568610
rect 90681 568568 90692 568582
rect 90748 568568 90759 568624
rect 90681 568566 90759 568568
rect 90969 566380 91047 566382
rect 90969 566366 90980 566380
rect 90590 566338 90980 566366
rect 90969 566324 90980 566338
rect 91036 566324 91047 566380
rect 90969 566322 91047 566324
rect 90767 564136 90845 564138
rect 90767 564122 90778 564136
rect 90586 564094 90778 564122
rect 90767 564080 90778 564094
rect 90834 564080 90845 564136
rect 90767 564078 90845 564080
rect 90757 561892 90835 561894
rect 90757 561878 90768 561892
rect 90590 561850 90768 561878
rect 90757 561836 90768 561850
rect 90824 561836 90835 561892
rect 90757 561834 90835 561836
rect 90715 559716 90793 559718
rect 90715 559702 90726 559716
rect 90588 559674 90726 559702
rect 90715 559660 90726 559674
rect 90782 559660 90793 559716
rect 90715 559658 90793 559660
rect 90739 557472 90817 557474
rect 90739 557458 90750 557472
rect 90590 557430 90750 557458
rect 90739 557416 90750 557430
rect 90806 557416 90817 557472
rect 90739 557414 90817 557416
rect 90673 555228 90751 555230
rect 90673 555214 90684 555228
rect 90588 555186 90684 555214
rect 90673 555172 90684 555186
rect 90740 555172 90751 555228
rect 90673 555170 90751 555172
rect 90707 552984 90785 552986
rect 90707 552970 90718 552984
rect 90586 552942 90718 552970
rect 90707 552928 90718 552942
rect 90774 552928 90785 552984
rect 90707 552926 90785 552928
rect 91840 550768 91952 587526
rect 93691 578391 93824 578421
rect 93691 578335 93729 578391
rect 93785 578335 93824 578391
rect 93691 578306 93824 578335
rect 74319 550726 74430 550768
rect 90754 550726 91952 550768
rect 74319 550698 74548 550726
rect 16692 468336 17076 468392
rect 17132 468336 17468 468392
rect 16692 468220 17468 468336
rect 22226 544230 23022 544294
rect 22226 544014 22562 544230
rect 22778 544014 23022 544230
rect 22226 425170 23022 544014
rect 29318 541794 29423 541808
rect 29312 541774 29423 541794
rect 29312 541718 29342 541774
rect 29398 541718 29423 541774
rect 29312 541685 29423 541718
rect 22226 425114 22644 425170
rect 22700 425114 23022 425170
rect 22226 425028 23022 425114
rect 26112 539466 27404 539534
rect 26112 539090 26546 539466
rect 26922 539090 27404 539466
rect 26112 295504 27404 539090
rect 29312 534306 29416 541685
rect 29303 534282 29425 534306
rect 29303 534226 29336 534282
rect 29392 534226 29425 534282
rect 29303 534202 29425 534226
rect 29312 530722 29416 534202
rect 74319 533152 74430 550698
rect 74734 550170 74762 550716
rect 74709 550168 74787 550170
rect 74709 550112 74720 550168
rect 74776 550112 74787 550168
rect 74709 550110 74787 550112
rect 82554 547470 82582 550718
rect 90374 550580 90402 550722
rect 90586 550698 91952 550726
rect 90754 550656 91952 550698
rect 82529 547468 82607 547470
rect 82529 547412 82540 547468
rect 82596 547412 82607 547468
rect 82529 547410 82607 547412
rect 90331 541804 90446 550580
rect 91840 544184 91952 550656
rect 91831 544156 91961 544184
rect 91831 544100 91868 544156
rect 91924 544100 91961 544156
rect 91831 544072 91961 544100
rect 90322 541774 90455 541804
rect 93700 541799 93815 578306
rect 101784 568092 101940 568111
rect 101784 567956 101794 568092
rect 101930 567956 101940 568092
rect 101363 566430 101521 566459
rect 101363 566294 101374 566430
rect 101510 566294 101521 566430
rect 100896 564180 101060 564203
rect 100896 564044 100910 564180
rect 101046 564044 101060 564180
rect 100463 561892 100593 561938
rect 100463 561836 100500 561892
rect 100556 561836 100593 561892
rect 99970 559692 100090 559733
rect 99970 559636 100002 559692
rect 100058 559636 100090 559692
rect 99470 557468 99598 557513
rect 99470 557412 99506 557468
rect 99562 557412 99598 557468
rect 99053 555230 99187 555278
rect 99053 555174 99092 555230
rect 99148 555174 99187 555230
rect 98621 552984 98755 553032
rect 98621 552928 98660 552984
rect 98716 552928 98755 552984
rect 90322 541718 90360 541774
rect 90416 541718 90455 541774
rect 90322 541689 90455 541718
rect 93696 541774 93819 541799
rect 93696 541718 93729 541774
rect 93785 541718 93819 541774
rect 93696 541694 93819 541718
rect 93700 541689 93815 541694
rect 74319 533096 74346 533152
rect 74402 533096 74430 533152
rect 74319 533060 74430 533096
rect 98621 532934 98755 552928
rect 98617 532900 98759 532934
rect 98617 532844 98660 532900
rect 98716 532844 98759 532900
rect 98617 532810 98759 532844
rect 98621 532805 98755 532810
rect 99053 532684 99187 555174
rect 99049 532650 99191 532684
rect 99049 532594 99092 532650
rect 99148 532594 99191 532650
rect 99049 532560 99191 532594
rect 99053 532555 99187 532560
rect 99470 532437 99598 557412
rect 99466 532406 99602 532437
rect 99466 532350 99506 532406
rect 99562 532350 99602 532406
rect 99466 532319 99602 532350
rect 99470 532314 99598 532319
rect 99970 532215 100090 559636
rect 99966 532188 100094 532215
rect 99966 532132 100002 532188
rect 100058 532132 100094 532188
rect 99966 532105 100094 532132
rect 99970 532100 100090 532105
rect 100463 531960 100593 561836
rect 100459 531928 100597 531960
rect 100459 531872 100500 531928
rect 100556 531872 100597 531928
rect 100459 531840 100597 531872
rect 100463 531835 100593 531840
rect 100896 531685 101060 564044
rect 100892 531676 101064 531685
rect 100892 531540 100910 531676
rect 101046 531540 101064 531676
rect 100892 531531 101064 531540
rect 100896 531526 101060 531531
rect 101363 531350 101521 566294
rect 101359 531344 101525 531350
rect 101359 531208 101374 531344
rect 101510 531208 101525 531344
rect 101359 531202 101525 531208
rect 101363 531197 101521 531202
rect 101784 531035 101940 567956
rect 183928 561633 184028 561638
rect 183924 561616 184032 561633
rect 183924 561560 183950 561616
rect 184006 561560 184032 561616
rect 183924 561543 184032 561560
rect 149940 556673 150040 556678
rect 149936 556656 150044 556673
rect 149936 556600 149962 556656
rect 150018 556600 150044 556656
rect 149936 556583 150044 556600
rect 149540 554689 149640 554694
rect 149536 554672 149644 554689
rect 149536 554616 149562 554672
rect 149618 554616 149644 554672
rect 149536 554599 149644 554616
rect 149540 549362 149640 554599
rect 149531 549340 149649 549362
rect 149531 549284 149562 549340
rect 149618 549284 149649 549340
rect 149531 549262 149649 549284
rect 149940 548618 150040 556583
rect 183928 555004 184028 561543
rect 251836 557534 251896 557543
rect 251836 557532 252104 557534
rect 251836 557476 251838 557532
rect 251894 557476 252104 557532
rect 251836 557474 252104 557476
rect 251836 557465 251896 557474
rect 226886 555249 227082 555254
rect 226882 555224 227086 555249
rect 226882 555088 226916 555224
rect 227052 555088 227086 555224
rect 226882 555063 227086 555088
rect 182912 554904 184028 555004
rect 182912 551026 183012 554904
rect 182903 551004 183021 551026
rect 182903 550948 182934 551004
rect 182990 550948 183021 551004
rect 182903 550926 183021 550948
rect 149931 548596 150049 548618
rect 225796 548612 225916 554692
rect 226886 552466 227082 555063
rect 226877 552436 227091 552466
rect 226877 552300 226916 552436
rect 227052 552300 227091 552436
rect 226877 552270 227091 552300
rect 323712 551121 324526 696231
rect 326095 693536 327363 693573
rect 326095 692360 326141 693536
rect 327317 692360 327363 693536
rect 326095 692323 327363 692360
rect 323712 550825 323936 551121
rect 324232 550825 324526 551121
rect 323712 550808 324526 550825
rect 326104 548756 327354 692323
rect 401679 691094 402065 699560
rect 417389 699226 417731 699258
rect 417389 698930 417412 699226
rect 417708 698930 417731 699226
rect 403319 697045 404123 697049
rect 414474 697045 415278 697049
rect 403314 697026 407485 697045
rect 403314 696250 403333 697026
rect 404109 696250 407485 697026
rect 403314 696231 407485 696250
rect 410401 697026 415283 697045
rect 410401 696250 414488 697026
rect 415264 696250 415283 697026
rect 410401 696231 415283 696250
rect 403319 696227 404123 696231
rect 414474 696227 415278 696231
rect 417389 693910 417731 698930
rect 470545 699226 470899 699264
rect 470545 698930 470574 699226
rect 470870 698930 470899 699226
rect 459850 696214 460194 696223
rect 459850 696190 461858 696214
rect 459850 695894 459874 696190
rect 460170 695894 461858 696190
rect 459850 695870 461858 695894
rect 459850 695861 460194 695870
rect 410642 693568 417731 693910
rect 467602 693328 468170 693337
rect 456947 693312 461852 693328
rect 456947 692776 456972 693312
rect 457508 692776 461852 693312
rect 456947 692760 461852 692776
rect 465516 693312 468170 693328
rect 465516 692776 467618 693312
rect 468154 692776 468170 693312
rect 465516 692760 468170 692776
rect 467602 692751 468170 692760
rect 401679 690718 401684 691094
rect 402060 690718 402065 691094
rect 401679 690622 402065 690718
rect 470545 690222 470899 698930
rect 562827 695682 574538 695684
rect 562827 695306 562838 695682
rect 563214 695306 574538 695682
rect 562827 695304 574538 695306
rect 569177 692878 569871 692882
rect 562085 692860 562779 692864
rect 562080 692816 564634 692860
rect 562080 692200 562124 692816
rect 562740 692200 564634 692816
rect 562080 692156 564634 692200
rect 567686 692834 569876 692878
rect 567686 692218 569216 692834
rect 569832 692218 569876 692834
rect 567686 692174 569876 692218
rect 569177 692170 569871 692174
rect 562085 692152 562779 692156
rect 465608 689868 470899 690222
rect 560028 689712 560392 689721
rect 560028 689678 571046 689712
rect 560028 689382 560062 689678
rect 560358 689382 571046 689678
rect 560028 689348 571046 689382
rect 560028 689339 560392 689348
rect 333289 683826 334011 683830
rect 333289 683130 333302 683826
rect 333998 683130 334011 683826
rect 333289 683126 334011 683130
rect 333298 632147 334002 683126
rect 570682 677644 571046 689348
rect 574158 683606 574538 695304
rect 574158 683226 575776 683606
rect 572977 680700 575276 680716
rect 572977 680164 573002 680700
rect 573538 680164 575276 680700
rect 572977 680148 575276 680164
rect 578940 680700 581133 680716
rect 578940 680164 580572 680700
rect 581108 680164 581133 680700
rect 578940 680148 581133 680164
rect 570682 677280 575342 677644
rect 567378 663569 567972 663581
rect 567378 663545 567987 663569
rect 567378 663009 567418 663545
rect 567954 663009 567987 663545
rect 567378 662985 567987 663009
rect 545434 633699 546234 633704
rect 545430 633692 546238 633699
rect 545430 632916 545446 633692
rect 546222 632916 546238 633692
rect 545430 632909 546238 632916
rect 333294 632108 334006 632147
rect 333294 631492 333342 632108
rect 333958 631492 334006 632108
rect 333294 631453 334006 631492
rect 333298 631448 334002 631453
rect 332399 627024 332909 627029
rect 332395 627002 332913 627024
rect 332395 626546 332426 627002
rect 332882 626546 332913 627002
rect 332395 626524 332913 626546
rect 330324 625953 331056 625958
rect 330320 625940 331060 625953
rect 330320 625244 330342 625940
rect 331038 625244 331060 625940
rect 330320 625231 331060 625244
rect 330324 618022 331056 625231
rect 330315 618004 331065 618022
rect 330315 617308 330342 618004
rect 331038 617308 331065 618004
rect 330315 617290 331065 617308
rect 332399 613019 332909 626524
rect 332390 612992 332918 613019
rect 332390 612536 332426 612992
rect 332882 612536 332918 612992
rect 332390 612509 332918 612536
rect 545434 582788 546234 632909
rect 545434 582012 545446 582788
rect 546222 582012 546234 582788
rect 545434 581991 546234 582012
rect 149931 548540 149962 548596
rect 150018 548540 150049 548596
rect 149931 548518 150049 548540
rect 225787 548580 225925 548612
rect 225787 548524 225828 548580
rect 225884 548524 225925 548580
rect 225787 548492 225925 548524
rect 326104 548300 326394 548756
rect 326850 548300 327354 548756
rect 326104 548212 327354 548300
rect 102435 547464 102583 547501
rect 102435 547408 102481 547464
rect 102537 547408 102583 547464
rect 102435 547371 102583 547408
rect 101780 531030 101944 531035
rect 101780 530894 101794 531030
rect 101930 530894 101944 531030
rect 102444 530990 102574 547371
rect 395919 536928 396051 536957
rect 395919 536872 395957 536928
rect 396013 536872 396051 536928
rect 395919 536843 396051 536872
rect 322595 535898 322755 535901
rect 322595 535762 322607 535898
rect 322743 535762 322755 535898
rect 322595 535759 322755 535762
rect 249181 534740 249317 534771
rect 249181 534684 249221 534740
rect 249277 534684 249317 534740
rect 249181 534653 249317 534684
rect 175851 533728 176009 533730
rect 175851 533592 175862 533728
rect 175998 533592 176009 533728
rect 175851 533590 176009 533592
rect 101780 530889 101944 530894
rect 101784 530884 101940 530889
rect 27853 530644 27931 530646
rect 27853 530588 27864 530644
rect 27920 530630 27931 530644
rect 27920 530602 29220 530630
rect 27920 530588 27931 530602
rect 27853 530586 27931 530588
rect 29350 530566 29378 530722
rect 102490 530568 102518 530990
rect 175860 530902 176000 533590
rect 175906 530560 175934 530902
rect 249190 530862 249308 534653
rect 322604 530890 322746 535759
rect 249230 530562 249258 530862
rect 322646 530560 322674 530890
rect 395928 530802 396042 536843
rect 542593 531464 542671 531466
rect 542593 531408 542604 531464
rect 542660 531408 542671 531464
rect 542593 531406 542671 531408
rect 469341 531043 469449 531060
rect 469341 530987 469367 531043
rect 469423 530987 469449 531043
rect 469341 530970 469449 530987
rect 395970 530562 395998 530802
rect 469350 530786 469440 530970
rect 469386 530564 469414 530786
rect 542618 530566 542646 531406
rect 552899 530658 552989 530667
rect 543074 530641 552989 530658
rect 543074 530630 552916 530641
rect 542772 530602 552916 530630
rect 543074 530585 552916 530602
rect 552972 530585 552989 530641
rect 543074 530568 552989 530585
rect 552899 530559 552989 530568
rect 27649 500452 27727 500454
rect 27649 500396 27660 500452
rect 27716 500438 27727 500452
rect 27716 500410 29214 500438
rect 27716 500396 27727 500410
rect 27649 500394 27727 500396
rect 27649 470260 27727 470262
rect 27649 470204 27660 470260
rect 27716 470246 27727 470260
rect 27716 470218 29214 470246
rect 27716 470204 27727 470218
rect 27649 470202 27727 470204
rect 27649 440068 27727 440070
rect 27649 440012 27660 440068
rect 27716 440054 27727 440068
rect 27716 440026 29214 440054
rect 27716 440012 27727 440026
rect 27649 440010 27727 440012
rect 27649 409944 27727 409946
rect 27649 409888 27660 409944
rect 27716 409930 27727 409944
rect 27716 409902 29214 409930
rect 27716 409888 27727 409902
rect 27649 409886 27727 409888
rect 27649 379752 27727 379754
rect 27649 379696 27660 379752
rect 27716 379738 27727 379752
rect 27716 379710 29214 379738
rect 27716 379696 27727 379710
rect 27649 379694 27727 379696
rect 27649 349560 27727 349562
rect 27649 349504 27660 349560
rect 27716 349546 27727 349560
rect 27716 349518 29214 349546
rect 27716 349504 27727 349518
rect 27649 349502 27727 349504
rect 27649 319436 27727 319438
rect 27649 319380 27660 319436
rect 27716 319422 27727 319436
rect 27716 319394 29214 319422
rect 27716 319380 27727 319394
rect 27649 319378 27727 319380
rect 26112 295448 26722 295504
rect 26778 295448 27404 295504
rect 26112 295414 27404 295448
rect 26586 289244 26646 289255
rect 26586 289188 26588 289244
rect 26644 289230 26646 289244
rect 26644 289202 29214 289230
rect 26644 289188 26646 289202
rect 26586 289177 26646 289188
rect 555728 274216 555788 274227
rect 555728 274202 555730 274216
rect 542778 274174 555730 274202
rect 555728 274160 555730 274174
rect 555786 274160 555788 274216
rect 555728 274149 555788 274160
rect 26818 259052 26878 259063
rect 26818 258996 26820 259052
rect 26876 259038 26878 259052
rect 26876 259010 29212 259038
rect 26876 258996 26878 259010
rect 26818 258985 26878 258996
rect 14310 248880 14626 248936
rect 14682 248880 14978 248936
rect 14310 248824 14978 248880
rect 27056 228860 27116 228871
rect 27056 228804 27058 228860
rect 27114 228846 27116 228860
rect 27114 228818 29220 228846
rect 27114 228804 27116 228818
rect 27056 228793 27116 228804
rect 27284 198736 27344 198747
rect 27284 198680 27286 198736
rect 27342 198722 27344 198736
rect 27342 198694 29214 198722
rect 27342 198680 27344 198694
rect 27284 198669 27344 198680
rect 27518 168544 27578 168555
rect 27518 168488 27520 168544
rect 27576 168530 27578 168544
rect 27576 168502 29212 168530
rect 27576 168488 27578 168502
rect 27518 168477 27578 168488
rect 27752 138352 27812 138363
rect 27752 138296 27754 138352
rect 27810 138338 27812 138352
rect 27810 138310 29210 138338
rect 27810 138296 27812 138310
rect 27752 138285 27812 138296
rect 9596 121258 10018 121314
rect 10074 121258 10498 121314
rect 9596 121187 10498 121258
rect 27976 108228 28036 108239
rect 27976 108172 27978 108228
rect 28034 108214 28036 108228
rect 28034 108186 29216 108214
rect 28034 108172 28036 108186
rect 27976 108161 28036 108172
rect 6634 81582 7188 81638
rect 7244 81582 7768 81638
rect 6634 81555 7768 81582
rect 28230 78036 28290 78047
rect 28230 77980 28232 78036
rect 28288 78022 28290 78036
rect 28288 77994 29214 78022
rect 28288 77980 28290 77994
rect 28230 77969 28290 77980
rect 567378 48180 567972 662985
rect 569844 662044 570372 662048
rect 569839 662003 580601 662044
rect 569839 661547 569880 662003
rect 570336 661547 580601 662003
rect 569839 661506 580601 661547
rect 569844 661502 570372 661506
rect 580063 92838 580601 661506
rect 580063 92782 580300 92838
rect 580356 92782 580601 92838
rect 580063 92707 580601 92782
rect 567378 48124 567626 48180
rect 567682 48124 567972 48180
rect 567378 48091 567972 48124
rect 28522 47844 28582 47855
rect 28522 47788 28524 47844
rect 28580 47830 28582 47844
rect 28580 47802 29220 47830
rect 28580 47788 28582 47802
rect 28522 47777 28582 47788
rect 28864 17720 28924 17731
rect 28864 17664 28866 17720
rect 28922 17706 28924 17720
rect 558978 17720 559038 17731
rect 558978 17706 558980 17720
rect 28922 17678 29230 17706
rect 542780 17678 558980 17706
rect 28922 17664 28924 17678
rect 28864 17653 28924 17664
rect 558978 17664 558980 17678
rect 559036 17664 559038 17720
rect 558978 17653 559038 17664
rect 579052 14662 579174 14668
rect 578190 14659 579174 14662
rect 578190 14629 579055 14659
rect 578190 14573 578232 14629
rect 578288 14573 579055 14629
rect 578190 14543 579055 14573
rect 579171 14543 579174 14659
rect 578190 14540 579174 14543
rect 578575 9936 578697 14540
rect 579052 14534 579174 14540
rect 580143 14659 580265 14668
rect 580143 14543 580146 14659
rect 580262 14658 580265 14659
rect 582049 14658 582151 14662
rect 580262 14630 582156 14658
rect 580262 14574 582072 14630
rect 582128 14574 582156 14630
rect 580262 14546 582156 14574
rect 580262 14543 580265 14546
rect 580143 14534 580265 14543
rect 582049 14542 582151 14546
rect 579064 9936 579186 9942
rect 578575 9933 579186 9936
rect 578575 9817 579067 9933
rect 579183 9817 579186 9933
rect 578575 9814 579186 9817
rect 578575 5206 578697 9814
rect 579064 9808 579186 9814
rect 580155 9933 580277 9942
rect 580155 9817 580158 9933
rect 580274 9932 580277 9933
rect 582061 9932 582163 9936
rect 580274 9904 582168 9932
rect 580274 9848 582084 9904
rect 582140 9848 582168 9904
rect 580274 9820 582168 9848
rect 580274 9817 580277 9820
rect 580155 9808 580277 9817
rect 582061 9816 582163 9820
rect 579176 5206 579298 5212
rect 578575 5203 579298 5206
rect 578575 5087 579179 5203
rect 579295 5087 579298 5203
rect 578575 5084 579298 5087
rect 578575 5075 578697 5084
rect 579176 5078 579298 5084
rect 580267 5203 580389 5212
rect 580267 5087 580270 5203
rect 580386 5202 580389 5203
rect 582173 5202 582275 5206
rect 580386 5174 582280 5202
rect 580386 5118 582196 5174
rect 582252 5118 582280 5174
rect 580386 5090 582280 5118
rect 580386 5087 580389 5090
rect 580267 5078 580389 5087
rect 582173 5086 582275 5090
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 171936 702024 171992 702080
rect 174442 702024 174498 702080
rect 223724 702024 223780 702080
rect 226124 702024 226180 702080
rect 325362 702024 325418 702080
rect 327872 702024 327928 702080
rect 26122 700224 26578 700680
rect 18332 697282 18708 697658
rect 28719 697242 29095 697618
rect 30210 694295 30586 694671
rect 9744 685562 10120 685938
rect 2923 682550 3219 682846
rect 9022 679578 9398 679954
rect 133206 698926 133502 699222
rect 122414 698444 122790 698820
rect 130768 698460 131144 698836
rect 70570 697302 70946 697678
rect 78990 697276 79366 697652
rect 82000 695454 82376 695830
rect 122502 695442 122798 695738
rect 71612 694279 71988 694655
rect 69202 690184 69578 690560
rect 171936 699052 171992 699108
rect 196563 700278 197099 700814
rect 174434 699054 174490 699110
rect 194114 697432 194570 697888
rect 186410 695070 186786 695446
rect 185248 694492 185384 694628
rect 134514 690190 134890 690566
rect 12334 679578 12710 679954
rect 4150 656518 5086 657454
rect 9619 658582 10475 659438
rect 7870 549135 8166 549431
rect 11780 654328 12636 655184
rect 9926 600492 10062 600628
rect 4626 338670 4682 338726
rect 7102 548396 7398 548692
rect 9980 547326 10196 547542
rect 90760 622094 90816 622150
rect 90676 619918 90732 619974
rect 90964 617674 91020 617730
rect 90762 615430 90818 615486
rect 90752 613186 90808 613242
rect 90710 611010 90766 611066
rect 90734 608766 90790 608822
rect 90668 606522 90724 606578
rect 90702 604278 90758 604334
rect 12260 381892 12316 381948
rect 14610 601188 14746 601324
rect 14590 550028 14806 550244
rect 16920 596647 17216 596943
rect 74704 601224 74760 601280
rect 98710 619912 98766 619968
rect 98396 617690 98452 617746
rect 98092 615434 98148 615490
rect 97788 613176 97844 613232
rect 97498 610968 97554 611024
rect 97218 608770 97274 608826
rect 96914 606514 96970 606570
rect 82524 600528 82580 600584
rect 74080 594474 74136 594530
rect 91852 596768 91908 596824
rect 96660 604280 96716 604336
rect 96660 594176 96716 594232
rect 96914 593880 96970 593936
rect 97218 593612 97274 593668
rect 97498 593342 97554 593398
rect 97788 593030 97844 593086
rect 98092 592740 98148 592796
rect 98396 592450 98452 592506
rect 185658 693166 185794 693302
rect 185288 617614 185344 617670
rect 219636 699858 220092 700314
rect 210686 695110 210982 695406
rect 221438 698926 221734 699222
rect 223720 699068 223776 699124
rect 264712 700324 264848 700460
rect 226118 699088 226174 699144
rect 209720 693592 210096 693968
rect 204982 692072 205278 692368
rect 202486 686483 202782 686779
rect 313095 700167 313711 700783
rect 321283 700174 321899 700790
rect 310840 698924 311136 699220
rect 314738 697578 315194 698034
rect 325370 699028 325426 699084
rect 327864 699040 327920 699096
rect 323731 696250 324507 697026
rect 282166 663222 282302 663358
rect 279761 661642 279817 661698
rect 215194 656798 215410 657014
rect 215904 654542 216120 654758
rect 222666 648334 222722 648390
rect 220316 638786 220372 638842
rect 220172 634256 220228 634312
rect 294494 640052 294550 640108
rect 285264 633934 285400 634070
rect 267210 632598 267346 632734
rect 244696 628530 244832 628666
rect 265774 628526 265910 628662
rect 285264 632310 285400 632446
rect 282638 631852 282694 631908
rect 289054 631852 289110 631908
rect 294068 629770 294284 629986
rect 292002 629398 292058 629454
rect 245703 628188 245839 628324
rect 267210 628188 267346 628324
rect 292002 626762 292058 626818
rect 294849 626546 295305 627002
rect 245732 625668 245788 625724
rect 294068 625524 294284 625740
rect 292242 623668 292298 623724
rect 294338 623668 294394 623724
rect 185698 617600 185754 617656
rect 186450 617406 186746 617702
rect 182750 615836 182806 615892
rect 183088 615430 183144 615486
rect 183088 607610 183144 607666
rect 182750 605626 182806 605682
rect 270596 595364 270652 595366
rect 270596 595312 270598 595364
rect 270598 595312 270650 595364
rect 270650 595312 270652 595364
rect 270596 595310 270652 595312
rect 98710 592180 98766 592236
rect 90346 578335 90402 578391
rect 90692 568568 90748 568624
rect 90980 566324 91036 566380
rect 90778 564080 90834 564136
rect 90768 561836 90824 561892
rect 90726 559660 90782 559716
rect 90750 557416 90806 557472
rect 90684 555172 90740 555228
rect 90718 552928 90774 552984
rect 93729 578335 93785 578391
rect 17076 468336 17132 468392
rect 22562 544014 22778 544230
rect 29342 541718 29398 541774
rect 22644 425114 22700 425170
rect 26546 539090 26922 539466
rect 29336 534226 29392 534282
rect 74720 550112 74776 550168
rect 82540 547412 82596 547468
rect 91868 544100 91924 544156
rect 101794 567956 101930 568092
rect 101374 566294 101510 566430
rect 100910 564044 101046 564180
rect 100500 561836 100556 561892
rect 100002 559636 100058 559692
rect 99506 557412 99562 557468
rect 99092 555174 99148 555230
rect 98660 552928 98716 552984
rect 90360 541718 90416 541774
rect 93729 541718 93785 541774
rect 74346 533096 74402 533152
rect 98660 532844 98716 532900
rect 99092 532594 99148 532650
rect 99506 532350 99562 532406
rect 100002 532132 100058 532188
rect 100500 531872 100556 531928
rect 100910 531540 101046 531676
rect 101374 531208 101510 531344
rect 183950 561560 184006 561616
rect 149962 556600 150018 556656
rect 149562 554616 149618 554672
rect 149562 549284 149618 549340
rect 251838 557476 251894 557532
rect 226916 555088 227052 555224
rect 182934 550948 182990 551004
rect 226916 552300 227052 552436
rect 326141 692360 327317 693536
rect 323936 550825 324232 551121
rect 417412 698930 417708 699226
rect 403333 696250 404109 697026
rect 414488 696250 415264 697026
rect 470574 698930 470870 699226
rect 459874 695894 460170 696190
rect 456972 692776 457508 693312
rect 467618 692776 468154 693312
rect 401684 690718 402060 691094
rect 562838 695306 563214 695682
rect 562124 692200 562740 692816
rect 569216 692218 569832 692834
rect 560062 689382 560358 689678
rect 333302 683130 333998 683826
rect 573002 680164 573538 680700
rect 580572 680164 581108 680700
rect 567418 663009 567954 663545
rect 545446 632916 546222 633692
rect 333342 631492 333958 632108
rect 332426 626546 332882 627002
rect 330342 625244 331038 625940
rect 330342 617308 331038 618004
rect 332426 612536 332882 612992
rect 545446 582012 546222 582788
rect 149962 548540 150018 548596
rect 225828 548524 225884 548580
rect 326394 548300 326850 548756
rect 102481 547408 102537 547464
rect 101794 530894 101930 531030
rect 395957 536872 396013 536928
rect 322607 535762 322743 535898
rect 249221 534684 249277 534740
rect 175862 533592 175998 533728
rect 27864 530588 27920 530644
rect 542604 531408 542660 531464
rect 469367 530987 469423 531043
rect 552916 530585 552972 530641
rect 27660 500396 27716 500452
rect 27660 470204 27716 470260
rect 27660 440012 27716 440068
rect 27660 409888 27716 409944
rect 27660 379696 27716 379752
rect 27660 349504 27716 349560
rect 27660 319380 27716 319436
rect 26722 295448 26778 295504
rect 26588 289188 26644 289244
rect 555730 274160 555786 274216
rect 26820 258996 26876 259052
rect 14626 248880 14682 248936
rect 27058 228804 27114 228860
rect 27286 198680 27342 198736
rect 27520 168488 27576 168544
rect 27754 138296 27810 138352
rect 10018 121258 10074 121314
rect 27978 108172 28034 108228
rect 7188 81582 7244 81638
rect 28232 77980 28288 78036
rect 569880 661547 570336 662003
rect 580300 92782 580356 92838
rect 567626 48124 567682 48180
rect 28524 47788 28580 47844
rect 28866 17664 28922 17720
rect 558980 17664 559036 17720
rect 578232 14573 578288 14629
rect 582072 14574 582128 14630
rect 582084 9848 582140 9904
rect 582196 5118 582252 5174
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 18305 697658 18735 702300
rect 26115 700680 26585 700687
rect 26115 700224 26122 700680
rect 26578 700224 26585 700680
rect 26115 700217 26585 700224
rect 18305 697282 18332 697658
rect 18708 697282 18735 697658
rect 18305 697255 18735 697282
rect 26120 691015 26580 700217
rect 70564 697678 70952 702300
rect 122372 698820 122832 702300
rect 167845 700837 168427 702300
rect 171820 702080 172132 702300
rect 171820 702024 171936 702080
rect 171992 702024 172132 702080
rect 171820 701948 172132 702024
rect 174326 702080 174638 702300
rect 174326 702024 174442 702080
rect 174498 702024 174638 702080
rect 174326 701948 174638 702024
rect 178141 700837 178723 702300
rect 196535 700837 197127 700842
rect 167845 700814 197127 700837
rect 167845 700278 196563 700814
rect 197099 700278 197127 700814
rect 219622 700340 220106 702300
rect 223608 702080 223920 702300
rect 223608 702024 223724 702080
rect 223780 702024 223920 702080
rect 223608 701948 223920 702024
rect 226008 702080 226320 702300
rect 226008 702024 226124 702080
rect 226180 702024 226320 702080
rect 226008 701948 226320 702024
rect 229792 700340 230276 702300
rect 321251 701312 321929 702300
rect 325246 702080 325558 702300
rect 325246 702024 325362 702080
rect 325418 702024 325558 702080
rect 325246 701948 325558 702024
rect 327756 702080 328068 702300
rect 327756 702024 327872 702080
rect 327928 702024 328068 702080
rect 327756 701948 328068 702024
rect 321254 700814 321929 701312
rect 331423 700814 332101 702300
rect 167845 700255 197127 700278
rect 196535 700250 197127 700255
rect 219588 700314 230276 700340
rect 219588 699872 219636 700314
rect 219622 699858 219636 699872
rect 220092 699872 230276 700314
rect 264508 700783 313742 700814
rect 264508 700460 313095 700783
rect 264508 700324 264712 700460
rect 264848 700324 313095 700460
rect 264508 700167 313095 700324
rect 313711 700167 313742 700783
rect 264508 700136 313742 700167
rect 321254 700790 332101 700814
rect 321254 700174 321283 700790
rect 321899 700174 332101 700790
rect 321254 700136 332101 700174
rect 220092 699858 220106 699872
rect 219622 699844 220106 699858
rect 220606 699856 230276 699872
rect 132958 699345 413253 699376
rect 132958 699222 412672 699345
rect 132958 698926 133206 699222
rect 133502 699110 221438 699222
rect 133502 699108 174434 699110
rect 133502 699052 171936 699108
rect 171992 699054 174434 699108
rect 174490 699054 221438 699110
rect 171992 699052 221438 699054
rect 133502 698926 221438 699052
rect 221734 699220 412672 699222
rect 221734 699144 310840 699220
rect 221734 699124 226118 699144
rect 221734 699068 223720 699124
rect 223776 699088 226118 699124
rect 226174 699088 310840 699144
rect 223776 699068 310840 699088
rect 221734 698926 310840 699068
rect 132958 698924 310840 698926
rect 311136 699096 412672 699220
rect 311136 699084 327864 699096
rect 311136 699028 325370 699084
rect 325426 699040 327864 699084
rect 327920 699040 412672 699096
rect 325426 699028 412672 699040
rect 311136 698924 412672 699028
rect 122372 698444 122414 698820
rect 122790 698444 122832 698820
rect 122372 698402 122832 698444
rect 130726 698836 131186 698878
rect 130726 698460 130768 698836
rect 131144 698460 131186 698836
rect 132958 698801 412672 698924
rect 413216 698801 413253 699345
rect 132958 698770 413253 698801
rect 28692 697618 29122 697665
rect 28692 697242 28719 697618
rect 29095 697242 29122 697618
rect 70564 697302 70570 697678
rect 70946 697302 70952 697678
rect 130726 697890 131186 698460
rect 314727 698034 315205 698045
rect 194107 697890 194577 697895
rect 130726 697888 194577 697890
rect 70564 697296 70952 697302
rect 78984 697652 79372 697658
rect 28692 693414 29122 697242
rect 78984 697276 78990 697652
rect 79366 697276 79372 697652
rect 130726 697432 194114 697888
rect 194570 697432 194577 697888
rect 314727 697578 314738 698034
rect 315194 697578 315205 698034
rect 314727 697567 315205 697578
rect 130726 697430 194577 697432
rect 194107 697425 194577 697430
rect 30008 694671 72188 694840
rect 30008 694295 30210 694671
rect 30586 694655 72188 694671
rect 30586 694295 71612 694655
rect 30008 694279 71612 694295
rect 71988 694279 72188 694655
rect 78984 694756 79372 697276
rect 81812 695830 122960 696102
rect 81812 695454 82000 695830
rect 82376 695738 122960 695830
rect 82376 695454 122502 695738
rect 81812 695442 122502 695454
rect 122798 695442 122960 695738
rect 81812 695194 122960 695442
rect 186403 695448 186793 695453
rect 186403 695446 211024 695448
rect 186403 695070 186410 695446
rect 186786 695406 211024 695446
rect 186786 695110 210686 695406
rect 210982 695110 211024 695406
rect 186786 695070 211024 695110
rect 186403 695068 211024 695070
rect 186403 695063 186793 695068
rect 78984 694628 185462 694756
rect 78984 694492 185248 694628
rect 185384 694492 185462 694628
rect 78984 694368 185462 694492
rect 30008 693984 72188 694279
rect 209709 693968 210107 693979
rect 209709 693592 209720 693968
rect 210096 693592 210107 693968
rect 209709 693581 210107 693592
rect 28692 693302 185918 693414
rect 28692 693166 185658 693302
rect 185794 693166 185918 693302
rect 28692 692984 185918 693166
rect 204957 692368 205303 692393
rect 204957 692072 204982 692368
rect 205278 692072 205303 692368
rect 67914 691015 183014 691032
rect 15173 690797 183014 691015
rect 15173 689933 30438 690797
rect 34822 690566 183014 690797
rect 34822 690560 134514 690566
rect 34822 690184 69202 690560
rect 69578 690190 134514 690560
rect 134890 690190 183014 690566
rect 69578 690184 183014 690190
rect 34822 689933 183014 690184
rect 15173 689748 183014 689933
rect 9727 685950 10137 685955
rect 15173 685950 16440 689748
rect 67914 689708 183014 689748
rect 9727 685938 16466 685950
rect 9727 685562 9744 685938
rect 10120 685562 16466 685938
rect 9727 685550 16466 685562
rect 9727 685545 10137 685550
rect -800 682855 1700 685242
rect 181690 683002 183014 689708
rect 202456 686804 202812 686809
rect 204957 686804 205303 692072
rect 209714 687274 210102 693581
rect 314732 687274 315200 697567
rect 323707 697045 324531 697050
rect 415421 697045 416235 702300
rect 417384 699235 417736 699260
rect 417384 698931 417408 699235
rect 417712 698931 417736 699235
rect 417384 698930 417412 698931
rect 417708 698930 417736 698931
rect 417384 698902 417736 698930
rect 323707 697026 404128 697045
rect 323707 696250 323731 697026
rect 324507 696250 403333 697026
rect 404109 696250 404128 697026
rect 323707 696231 404128 696250
rect 414450 697026 416235 697045
rect 414450 696250 414488 697026
rect 415264 696250 416235 697026
rect 414450 696231 416235 696250
rect 323707 696226 324531 696231
rect 459845 696190 460199 696219
rect 459845 695894 459874 696190
rect 460170 695894 460199 696190
rect 459845 695865 460199 695894
rect 326099 693573 327359 693578
rect 326099 693536 457696 693573
rect 326099 692360 326141 693536
rect 327317 693312 457696 693536
rect 327317 692776 456972 693312
rect 457508 692776 457696 693312
rect 327317 692360 457696 692776
rect 326099 692323 457696 692360
rect 326099 692318 327359 692323
rect 401674 691094 402070 691104
rect 401674 690718 401684 691094
rect 402060 690718 402070 691094
rect 401674 690708 402070 690718
rect 401679 687274 402065 690708
rect 459850 687274 460194 695865
rect 467273 693312 468523 702300
rect 470540 699235 470904 699266
rect 470540 698931 470570 699235
rect 470874 698931 470904 699235
rect 470540 698930 470574 698931
rect 470870 698930 470904 698931
rect 470540 698896 470904 698930
rect 512816 699204 515276 702340
rect 520594 699204 523054 702340
rect 566594 702300 571594 704800
rect 512816 699166 523054 699204
rect 467273 692776 467618 693312
rect 468154 692776 468523 693312
rect 467273 692705 468523 692776
rect 512816 696782 520606 699166
rect 522990 696782 523054 699166
rect 512816 696744 523054 696782
rect 512816 695048 515276 696744
rect 512816 692664 512854 695048
rect 515238 692664 515276 695048
rect 512816 692620 515276 692664
rect 555818 695682 563468 696048
rect 555818 695306 562838 695682
rect 563214 695306 563468 695682
rect 555818 694724 563468 695306
rect 555818 687274 557142 694724
rect 562080 692816 562784 692860
rect 562080 692200 562124 692816
rect 562740 692200 562784 692816
rect 560023 689687 560397 689723
rect 560023 689383 560058 689687
rect 560362 689383 560397 689687
rect 560023 689382 560062 689383
rect 560358 689382 560397 689383
rect 560023 689343 560397 689382
rect 202456 686779 205303 686804
rect 202456 686483 202486 686779
rect 202782 686483 205303 686779
rect 202456 686458 205303 686483
rect 202456 686453 202812 686458
rect 207618 685950 557142 687274
rect 207618 683002 208942 685950
rect 333293 683830 334007 683835
rect 562080 683830 562784 692200
rect 569172 692834 569876 702300
rect 569172 692218 569216 692834
rect 569832 692218 569876 692834
rect 569172 692174 569876 692218
rect 333293 683826 562784 683830
rect 333293 683130 333302 683826
rect 333998 683130 562784 683826
rect 333293 683126 562784 683130
rect 333293 683121 334007 683126
rect -800 682846 3228 682855
rect -800 682550 2923 682846
rect 3219 682550 3228 682846
rect -800 682541 3228 682550
rect -800 680242 1700 682541
rect 181690 681678 208942 683002
rect 582300 680761 584800 682984
rect 572285 680700 573670 680761
rect 572285 680164 573002 680700
rect 573538 680164 573670 680700
rect 572285 680039 573670 680164
rect 580494 680700 584800 680761
rect 580494 680164 580572 680700
rect 581108 680164 584800 680700
rect 580494 680039 584800 680164
rect 12312 679971 12732 679976
rect 9005 679954 12732 679971
rect 9005 679578 9022 679954
rect 9398 679578 12334 679954
rect 12710 679578 12732 679954
rect 9005 679561 12732 679578
rect 12312 679556 12732 679561
rect 282128 663545 567983 663574
rect 282128 663358 567418 663545
rect 282128 663222 282166 663358
rect 282302 663222 567418 663358
rect 282128 663009 567418 663222
rect 567954 663009 567983 663545
rect 282128 662980 567983 663009
rect 279734 662003 570377 662044
rect 279734 661698 569880 662003
rect 279734 661642 279761 661698
rect 279817 661642 569880 661698
rect 279734 661547 569880 661642
rect 570336 661547 570377 662003
rect 279734 661506 570377 661547
rect 9475 659438 222804 659540
rect 9475 658582 9619 659438
rect 10475 658582 222804 659438
rect 9475 658398 222804 658582
rect 4122 657454 215506 657482
rect 4122 656518 4150 657454
rect 5086 657014 215506 657454
rect 5086 656798 215194 657014
rect 215410 656798 215506 657014
rect 5086 656518 215506 656798
rect 4122 656490 215506 656518
rect 11758 655184 216158 655206
rect 11758 654328 11780 655184
rect 12636 654758 216158 655184
rect 12636 654542 215904 654758
rect 216120 654542 216158 654758
rect 12636 654328 216158 654542
rect 11758 654306 216158 654328
rect -800 648564 1660 648642
rect -800 648544 19672 648564
rect -800 643920 15022 648544
rect 19646 643920 19672 648544
rect 222572 648390 222802 658398
rect 222572 648334 222666 648390
rect 222722 648334 222802 648390
rect 222572 648260 222802 648334
rect -800 643900 19672 643920
rect -800 643842 1660 643900
rect -800 638558 1660 638642
rect 8408 638558 13072 643900
rect 294472 640108 297043 640136
rect 294472 640052 294494 640108
rect 294550 640052 297043 640108
rect 294472 639998 297043 640052
rect 220294 638842 220600 638864
rect 220294 638786 220316 638842
rect 220372 638786 220600 638842
rect 220294 638764 220600 638786
rect -800 633894 13072 638558
rect 220150 634312 220420 634334
rect 220150 634256 220172 634312
rect 220228 634256 220420 634312
rect 220150 634234 220420 634256
rect 281465 634070 285433 634103
rect 281465 633934 285264 634070
rect 285400 633934 285433 634070
rect 281465 633901 285433 633934
rect -800 633842 1660 633894
rect 267172 632767 267384 632772
rect 281465 632767 281667 633901
rect 296905 633393 297043 639998
rect 321650 633692 546234 633704
rect 321650 633393 545446 633692
rect 296905 633255 545446 633393
rect 321650 632916 545446 633255
rect 546222 632916 546234 633692
rect 321650 632904 546234 632916
rect 267172 632734 281667 632767
rect 267172 632598 267210 632734
rect 267346 632598 281667 632734
rect 267172 632565 281667 632598
rect 267172 632560 267384 632565
rect 285226 632479 285438 632484
rect 285226 632446 289887 632479
rect 285226 632310 285264 632446
rect 285400 632310 289887 632446
rect 285226 632277 289887 632310
rect 285226 632272 285438 632277
rect 282611 631930 282721 631935
rect 282611 631908 289132 631930
rect 282611 631852 282638 631908
rect 282694 631852 289054 631908
rect 289110 631852 289132 631908
rect 282611 631830 289132 631852
rect 289685 631921 289887 632277
rect 329060 632108 334076 632152
rect 329060 631921 333342 632108
rect 282611 631825 282721 631830
rect 289685 631719 333342 631921
rect 270312 631406 289469 631592
rect 329060 631492 333342 631719
rect 333958 631492 334076 632108
rect 329060 631448 334076 631492
rect 270314 628860 270414 631406
rect 289283 630453 289469 631406
rect 572285 630692 573007 680039
rect 582300 677984 584800 680039
rect 582340 644550 584800 644584
rect 575932 644542 584800 644550
rect 575932 639838 575946 644542
rect 580650 639838 584800 644542
rect 575932 639830 584800 639838
rect 328964 630453 573007 630692
rect 577382 632996 579842 639830
rect 582340 639784 584800 639830
rect 582340 632996 584800 634584
rect 577382 630536 584800 632996
rect 289283 630267 573007 630453
rect 292322 629986 294304 630006
rect 292322 629928 294068 629986
rect 288724 629828 294068 629928
rect 292322 629770 294068 629828
rect 294284 629770 294304 629986
rect 328964 629970 573007 630267
rect 582340 629784 584800 630536
rect 292322 629750 294304 629770
rect 291952 629454 328227 629556
rect 291952 629398 292002 629454
rect 292058 629398 328227 629454
rect 291952 629310 328227 629398
rect 244667 628690 244861 628695
rect 265745 628690 265939 628691
rect 244667 628666 265950 628690
rect 244667 628530 244696 628666
rect 244832 628662 265950 628666
rect 244832 628530 265774 628662
rect 244667 628526 265774 628530
rect 265910 628526 265950 628662
rect 244667 628506 265950 628526
rect 244667 628501 244861 628506
rect 265745 628497 265939 628506
rect 327981 628382 328227 629310
rect 245665 628357 245877 628362
rect 245665 628324 267379 628357
rect 245665 628188 245703 628324
rect 245839 628188 267210 628324
rect 267346 628188 267379 628324
rect 245665 628155 267379 628188
rect 245665 628150 245877 628155
rect 327981 627637 577818 628382
rect 328008 627634 577818 627637
rect 294817 627029 295337 627034
rect 294817 627002 332909 627029
rect 268576 626818 292080 626840
rect 268576 626762 292002 626818
rect 292058 626762 292080 626818
rect 268576 626740 292080 626762
rect 294817 626546 294849 627002
rect 295305 626546 332426 627002
rect 332882 626546 332909 627002
rect 294817 626519 332909 626546
rect 294817 626514 295337 626519
rect 294006 625940 331056 625958
rect 245710 625724 245810 625746
rect 245710 625668 245732 625724
rect 245788 625668 245810 625724
rect 245710 625646 245810 625668
rect 294006 625740 330342 625940
rect 294006 625524 294068 625740
rect 294284 625524 330342 625740
rect 294006 625244 330342 625524
rect 331038 625244 331056 625940
rect 294006 625226 331056 625244
rect 292048 623724 292320 623746
rect 292048 623668 292242 623724
rect 292298 623668 292320 623724
rect 292048 623646 292320 623668
rect 294290 623724 574212 623952
rect 294290 623668 294338 623724
rect 294394 623668 574212 623724
rect 294290 623396 574212 623668
rect 90730 622150 93205 622204
rect 90730 622094 90760 622150
rect 90816 622094 93205 622150
rect 90730 622054 93205 622094
rect 93055 620431 93205 622054
rect 292480 621874 292580 623004
rect 292476 621228 569437 621874
rect 93055 620428 137997 620431
rect 93055 620284 137844 620428
rect 137988 620284 137997 620428
rect 93055 620281 137997 620284
rect 140292 620428 140440 620436
rect 140292 620284 140294 620428
rect 140438 620284 140440 620428
rect 140292 620276 140440 620284
rect 90649 619974 137091 620037
rect 90649 619918 90676 619974
rect 90732 619968 137091 619974
rect 90732 619918 98710 619968
rect 90649 619912 98710 619918
rect 98766 619912 137091 619968
rect 90649 619859 137091 619912
rect 90925 617746 135727 617803
rect 90925 617730 98396 617746
rect 90925 617674 90964 617730
rect 91020 617690 98396 617730
rect 98452 617690 135727 617746
rect 91020 617674 135727 617690
rect 90925 617625 135727 617674
rect 90737 615490 134349 615543
rect 90737 615486 98092 615490
rect 90737 615430 90762 615486
rect 90818 615434 98092 615486
rect 98148 615434 134349 615490
rect 90818 615430 134349 615434
rect 90737 615365 134349 615430
rect 90723 613242 132889 613299
rect 90723 613186 90752 613242
rect 90808 613232 132889 613242
rect 90808 613186 97788 613232
rect 90723 613176 97788 613186
rect 97844 613176 132889 613232
rect 90723 613121 132889 613176
rect 90679 611066 131559 611103
rect 90679 611010 90710 611066
rect 90766 611024 131559 611066
rect 90766 611010 97498 611024
rect 90679 610968 97498 611010
rect 97554 610968 131559 611024
rect 90679 610925 131559 610968
rect 90707 608826 130513 608885
rect 90707 608822 97218 608826
rect 90707 608766 90734 608822
rect 90790 608770 97218 608822
rect 97274 608770 130513 608826
rect 90790 608766 130513 608770
rect 90707 608707 130513 608766
rect 90647 606600 129595 606637
rect 90646 606578 129595 606600
rect 90646 606522 90668 606578
rect 90724 606570 129595 606578
rect 90724 606522 96914 606570
rect 90646 606514 96914 606522
rect 96970 606514 129595 606570
rect 90646 606504 129595 606514
rect 90647 606459 129595 606504
rect 90677 604336 128845 604395
rect 90677 604334 96660 604336
rect 90677 604278 90702 604334
rect 90758 604280 96660 604334
rect 96716 604280 128845 604336
rect 90758 604278 128845 604280
rect 90677 604217 128845 604278
rect 128667 602614 128845 604217
rect 129417 602912 129595 606459
rect 130335 603190 130513 608707
rect 131381 603472 131559 610925
rect 132711 603774 132889 613121
rect 134171 604048 134349 615365
rect 135549 604364 135727 617625
rect 136913 604652 137091 619859
rect 330319 618022 331061 618027
rect 330319 618004 563858 618022
rect 186408 617702 186788 617744
rect 185266 617670 185366 617692
rect 185266 617614 185288 617670
rect 185344 617614 185366 617670
rect 182723 615914 182833 615919
rect 185266 615914 185366 617614
rect 182723 615892 185366 615914
rect 182723 615836 182750 615892
rect 182806 615836 185366 615892
rect 182723 615814 185366 615836
rect 185676 617656 185776 617678
rect 185676 617600 185698 617656
rect 185754 617600 185776 617656
rect 182723 615809 182833 615814
rect 183061 615508 183171 615513
rect 185676 615508 185776 617600
rect 183061 615486 185776 615508
rect 183061 615430 183088 615486
rect 183144 615430 185776 615486
rect 183061 615408 185776 615430
rect 186408 617406 186450 617702
rect 186746 617406 186788 617702
rect 183061 615403 183171 615408
rect 186408 612782 186788 617406
rect 330319 617308 330342 618004
rect 331038 617308 563858 618004
rect 330319 617290 563858 617308
rect 330319 617285 331061 617290
rect 181778 612402 186788 612782
rect 332352 612992 558426 613476
rect 332352 612536 332426 612992
rect 332882 612536 558426 612992
rect 332352 611640 558426 612536
rect 181472 607666 183166 607688
rect 181472 607610 183088 607666
rect 183144 607610 183166 607666
rect 181472 607588 183166 607610
rect 181192 605682 182828 605704
rect 181192 605626 182750 605682
rect 182806 605626 182828 605682
rect 181192 605604 182828 605626
rect 136913 604474 142902 604652
rect 135549 604186 142904 604364
rect 134171 603870 142912 604048
rect 132711 603596 142914 603774
rect 131381 603294 142898 603472
rect 130335 603012 142894 603190
rect 129417 602734 142912 602912
rect 128667 602436 142914 602614
rect 14570 601324 74802 601364
rect 14570 601188 14610 601324
rect 14746 601280 74802 601324
rect 14746 601224 74704 601280
rect 74760 601224 74802 601280
rect 14746 601188 74802 601224
rect 14570 601148 74802 601188
rect 9890 600628 82612 600664
rect 9890 600492 9926 600628
rect 10062 600584 82612 600628
rect 10062 600528 82524 600584
rect 82580 600528 82612 600584
rect 10062 600492 82612 600528
rect 9890 600456 82612 600492
rect 16893 596943 91972 596970
rect 16893 596647 16920 596943
rect 17216 596824 91972 596943
rect 17216 596768 91852 596824
rect 91908 596768 91972 596824
rect 17216 596647 91972 596768
rect 16893 596620 91972 596647
rect 270283 595366 270674 595388
rect 270283 595310 270596 595366
rect 270652 595310 270674 595366
rect 270283 595288 270674 595310
rect 24254 594565 24386 594570
rect 74045 594565 74172 594566
rect 24253 594530 74179 594565
rect 24253 594466 24288 594530
rect 24352 594474 74080 594530
rect 74136 594474 74179 594530
rect 24352 594466 74179 594474
rect 24253 594431 74179 594466
rect 24254 594426 24386 594431
rect 24594 594263 24710 594268
rect 24593 594236 96747 594263
rect 24593 594172 24620 594236
rect 24684 594232 96747 594236
rect 24684 594176 96660 594232
rect 96716 594176 96747 594232
rect 24684 594172 96747 594176
rect 24593 594145 96747 594172
rect 24594 594140 24710 594145
rect 24914 593967 25030 593972
rect 24913 593940 97001 593967
rect 24913 593876 24940 593940
rect 25004 593936 97001 593940
rect 25004 593880 96914 593936
rect 96970 593880 97001 593936
rect 25004 593876 97001 593880
rect 24913 593849 97001 593876
rect 24914 593844 25030 593849
rect 25216 593699 25332 593704
rect 25215 593672 97305 593699
rect 25215 593608 25242 593672
rect 25306 593668 97305 593672
rect 25306 593612 97218 593668
rect 97274 593612 97305 593668
rect 25306 593608 97305 593612
rect 25215 593581 97305 593608
rect 25216 593576 25332 593581
rect 25494 593429 25610 593434
rect 25493 593402 97585 593429
rect 25493 593338 25520 593402
rect 25584 593398 97585 593402
rect 25584 593342 97498 593398
rect 97554 593342 97585 593398
rect 25584 593338 97585 593342
rect 25493 593311 97585 593338
rect 25494 593306 25610 593311
rect 25784 593117 25900 593122
rect 25783 593090 97875 593117
rect 25783 593026 25810 593090
rect 25874 593086 97875 593090
rect 25874 593030 97788 593086
rect 97844 593030 97875 593086
rect 25874 593026 97875 593030
rect 25783 592999 97875 593026
rect 25784 592994 25900 592999
rect 26066 592827 26182 592832
rect 26065 592800 98179 592827
rect 26065 592736 26092 592800
rect 26156 592796 98179 592800
rect 26156 592740 98092 592796
rect 98148 592740 98179 592796
rect 26156 592736 98179 592740
rect 26065 592709 98179 592736
rect 26066 592704 26182 592709
rect 26318 592537 26434 592542
rect 26317 592510 98483 592537
rect 26317 592446 26344 592510
rect 26408 592506 98483 592510
rect 26408 592450 98396 592506
rect 98452 592450 98483 592506
rect 26408 592446 98483 592450
rect 26317 592419 98483 592446
rect 26318 592414 26434 592419
rect 26555 592268 26673 592273
rect 26554 592240 98798 592268
rect 26554 592176 26582 592240
rect 26646 592236 98798 592240
rect 26646 592180 98710 592236
rect 98766 592180 98798 592236
rect 26646 592176 98798 592180
rect 26554 592148 98798 592176
rect 26555 592143 26673 592148
rect 270283 588060 270478 595288
rect 270282 588052 548702 588060
rect 270282 587608 552174 588052
rect 544900 582788 547088 582992
rect 544900 582012 545446 582788
rect 546222 582012 547088 582788
rect 93695 578421 93820 578426
rect 90317 578391 93820 578421
rect 90317 578335 90346 578391
rect 90402 578335 93729 578391
rect 93785 578335 93820 578391
rect 90317 578306 93820 578335
rect 93695 578301 93820 578306
rect 90651 568624 90928 568687
rect 90651 568568 90692 568624
rect 90748 568568 90928 568624
rect 90651 568509 90928 568568
rect 90750 568121 90928 568509
rect 90750 568092 137107 568121
rect 90750 567956 101794 568092
rect 101930 567956 137107 568092
rect 90750 567943 137107 567956
rect 101779 567941 101945 567943
rect 90941 566430 135743 566453
rect 90941 566380 101374 566430
rect 90941 566324 90980 566380
rect 91036 566324 101374 566380
rect 90941 566294 101374 566324
rect 101510 566294 135743 566430
rect 90941 566275 135743 566294
rect -800 559442 1660 564242
rect 100891 564193 101065 564199
rect 90753 564180 134365 564193
rect 90753 564136 100910 564180
rect 90753 564080 90778 564136
rect 90834 564080 100910 564136
rect 90753 564044 100910 564080
rect 101046 564044 134365 564180
rect 90753 564015 134365 564044
rect 90739 561892 132905 561949
rect 90739 561836 90768 561892
rect 90824 561836 100500 561892
rect 100556 561836 132905 561892
rect 90739 561771 132905 561836
rect 90695 559716 131575 559753
rect 90695 559660 90726 559716
rect 90782 559692 131575 559716
rect 90782 559660 100002 559692
rect 90695 559636 100002 559660
rect 100058 559636 131575 559692
rect 90695 559575 131575 559636
rect 90723 557525 99459 557535
rect 99742 557525 130529 557535
rect 90723 557472 130529 557525
rect 90723 557416 90750 557472
rect 90806 557468 130529 557472
rect 90806 557416 99506 557468
rect 90723 557412 99506 557416
rect 99562 557412 130529 557468
rect 90723 557366 130529 557412
rect 90723 557357 99459 557366
rect 99742 557357 130529 557366
rect 90663 555250 129611 555287
rect 90662 555230 129611 555250
rect 90662 555228 99092 555230
rect 90662 555172 90684 555228
rect 90740 555174 99092 555228
rect 99148 555174 129611 555230
rect 90740 555172 129611 555174
rect 90662 555154 129611 555172
rect 90663 555109 129611 555154
rect -800 549442 1660 554242
rect 90693 552984 128861 553045
rect 90693 552928 90718 552984
rect 90774 552928 98660 552984
rect 98716 552928 128861 552984
rect 90693 552867 128861 552928
rect 128683 551264 128861 552867
rect 129433 551562 129611 555109
rect 130351 551840 130529 557357
rect 131397 552122 131575 559575
rect 132727 552424 132905 561771
rect 134187 552698 134365 564015
rect 135565 553014 135743 566275
rect 136929 553302 137107 567943
rect 183928 561616 184028 561832
rect 183928 561560 183950 561616
rect 184006 561560 184028 561616
rect 183928 561538 184028 561560
rect 251770 557532 251966 557566
rect 251770 557476 251838 557532
rect 251894 557476 251966 557532
rect 149940 556656 150040 556678
rect 149940 556600 149962 556656
rect 150018 556600 150040 556656
rect 149940 556578 150040 556600
rect 226886 555852 250874 556048
rect 226886 555224 227082 555852
rect 250678 555744 250874 555852
rect 251770 555744 251966 557476
rect 250678 555548 251966 555744
rect 226886 555088 226916 555224
rect 227052 555088 227082 555224
rect 226886 555058 227082 555088
rect 149540 554672 149640 554694
rect 149540 554616 149562 554672
rect 149618 554616 149640 554672
rect 149540 554594 149640 554616
rect 136929 553124 142918 553302
rect 142360 553122 142906 553124
rect 135565 552836 142920 553014
rect 142362 552834 142908 552836
rect 134187 552520 142928 552698
rect 142370 552518 142916 552520
rect 180682 552436 227148 552576
rect 132727 552246 142930 552424
rect 180682 552300 226916 552436
rect 227052 552300 227148 552436
rect 142372 552244 142918 552246
rect 131397 551944 142914 552122
rect 180682 552120 227148 552300
rect 142356 551942 142902 551944
rect 130351 551662 142910 551840
rect 142352 551660 142898 551662
rect 129433 551384 142928 551562
rect 142370 551382 142916 551384
rect 128683 551086 142930 551264
rect 142372 551084 142918 551086
rect 14568 550244 74810 550266
rect 14568 550028 14590 550244
rect 14806 550168 74810 550244
rect 14806 550112 74720 550168
rect 74776 550112 74810 550168
rect 14806 550028 74810 550112
rect 14568 550006 74810 550028
rect 7861 549431 149688 549440
rect 7861 549135 7870 549431
rect 8166 549340 149688 549431
rect 8166 549284 149562 549340
rect 149618 549284 149688 549340
rect 8166 549135 149688 549284
rect 7861 549126 149688 549135
rect 7074 548692 150086 548720
rect 7074 548396 7102 548692
rect 7398 548596 150086 548692
rect 7398 548540 149962 548596
rect 150018 548540 150086 548596
rect 7398 548396 150086 548540
rect 7074 548368 150086 548396
rect 9958 547542 102608 547564
rect 9958 547326 9980 547542
rect 10196 547468 102608 547542
rect 10196 547412 82540 547468
rect 82596 547464 102608 547468
rect 82596 547412 102481 547464
rect 10196 547408 102481 547412
rect 102537 547408 102608 547464
rect 10196 547326 102608 547408
rect 9958 547304 102608 547326
rect 22538 544230 92000 544254
rect 22538 544014 22562 544230
rect 22778 544156 92000 544230
rect 22778 544100 91868 544156
rect 91924 544100 92000 544156
rect 22778 544014 92000 544100
rect 22538 543990 92000 544014
rect 90326 541804 90451 541809
rect 29313 541774 93815 541804
rect 29313 541718 29342 541774
rect 29398 541718 90360 541774
rect 90416 541718 93729 541774
rect 93785 541718 93815 541774
rect 29313 541689 93815 541718
rect 90326 541684 90451 541689
rect 180682 539506 181138 552120
rect 182880 551121 324243 551132
rect 182880 551004 323936 551121
rect 182880 550948 182934 551004
rect 182990 550948 323936 551004
rect 182880 550825 323936 550948
rect 324232 550825 324243 551121
rect 182880 550814 324243 550825
rect 225694 548756 326874 548780
rect 225694 548580 326394 548756
rect 225694 548524 225828 548580
rect 225884 548524 326394 548580
rect 225694 548300 326394 548524
rect 326850 548300 326874 548756
rect 225694 548276 326874 548300
rect 26506 539466 181138 539506
rect 26506 539090 26546 539466
rect 26922 539090 181138 539466
rect 26506 539050 181138 539090
rect 20195 537048 20473 537054
rect 20195 537021 396092 537048
rect 20195 536797 20222 537021
rect 20446 536928 396092 537021
rect 20446 536872 395957 536928
rect 396013 536872 396092 536928
rect 20446 536797 396092 536872
rect 20195 536770 396092 536797
rect 20195 536764 20473 536770
rect 21652 536092 22172 536098
rect 21652 536064 322800 536092
rect 21652 535600 21680 536064
rect 22144 535898 322800 536064
rect 22144 535762 322607 535898
rect 322743 535762 322800 535898
rect 22144 535600 322800 535762
rect 21652 535572 322800 535600
rect 21652 535566 22172 535572
rect 22676 534894 23016 534900
rect 22676 534876 249362 534894
rect 22676 534572 22694 534876
rect 22998 534740 249362 534876
rect 22998 534684 249221 534740
rect 249277 534684 249362 534740
rect 22998 534572 249362 534684
rect 22676 534554 249362 534572
rect 22676 534548 23016 534554
rect 29307 534306 29421 534311
rect 19726 534282 29421 534306
rect 19726 534226 29336 534282
rect 29392 534226 29421 534282
rect 19726 534202 29421 534226
rect -800 511530 484 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect 19726 508096 19830 534202
rect 29307 534197 29421 534202
rect 23489 533848 23855 533854
rect 23489 533817 176034 533848
rect 23489 533513 23520 533817
rect 23824 533728 176034 533817
rect 23824 533592 175862 533728
rect 175998 533592 176034 533728
rect 23824 533513 176034 533592
rect 23489 533482 176034 533513
rect 23489 533476 23855 533482
rect 26785 533179 26913 533184
rect 74314 533179 74435 533185
rect 26784 533152 74455 533179
rect 26784 533146 74346 533152
rect 26784 533082 26817 533146
rect 26881 533096 74346 533146
rect 74402 533096 74455 533152
rect 26881 533082 74455 533096
rect 26784 533049 74455 533082
rect 26785 533044 26913 533049
rect 27019 532939 27151 532944
rect 27018 532904 98755 532939
rect 27018 532840 27053 532904
rect 27117 532900 98755 532904
rect 27117 532844 98660 532900
rect 98716 532844 98755 532900
rect 27117 532840 98755 532844
rect 27018 532805 98755 532840
rect 27019 532800 27151 532805
rect 27247 532689 27379 532694
rect 27246 532654 99187 532689
rect 27246 532590 27281 532654
rect 27345 532650 99187 532654
rect 27345 532594 99092 532650
rect 99148 532594 99187 532650
rect 27345 532590 99187 532594
rect 27246 532555 99187 532590
rect 27247 532550 27379 532555
rect 27483 532442 27609 532447
rect 27482 532410 99598 532442
rect 27482 532346 27514 532410
rect 27578 532406 99598 532410
rect 27578 532350 99506 532406
rect 99562 532350 99598 532406
rect 27578 532346 99598 532350
rect 27482 532314 99598 532346
rect 27483 532309 27609 532314
rect 27715 532220 27833 532225
rect 27714 532192 100090 532220
rect 27714 532128 27742 532192
rect 27806 532188 100090 532192
rect 27806 532132 100002 532188
rect 100058 532132 100090 532188
rect 27806 532128 100090 532132
rect 27714 532100 100090 532128
rect 27715 532095 27833 532100
rect 27945 531965 28073 531970
rect 27944 531932 100593 531965
rect 27944 531868 27977 531932
rect 28041 531928 100593 531932
rect 28041 531872 100500 531928
rect 100556 531872 100593 531928
rect 28041 531868 100593 531872
rect 27944 531835 100593 531868
rect 27945 531830 28073 531835
rect 28177 531690 28339 531695
rect 28176 531680 101060 531690
rect 28176 531536 28186 531680
rect 28330 531676 101060 531680
rect 28330 531540 100910 531676
rect 101046 531540 101060 531676
rect 28330 531536 101060 531540
rect 28176 531526 101060 531536
rect 28177 531521 28339 531526
rect 542574 531509 543627 531538
rect 542574 531464 543448 531509
rect 542574 531408 542604 531464
rect 542660 531408 543448 531464
rect 542574 531365 543448 531408
rect 543592 531365 543627 531509
rect 28483 531355 28639 531360
rect 28482 531348 101521 531355
rect 28482 531204 28489 531348
rect 28633 531344 101521 531348
rect 28633 531208 101374 531344
rect 101510 531208 101521 531344
rect 542574 531336 543627 531365
rect 28633 531204 101521 531208
rect 28482 531197 101521 531204
rect 28483 531192 28639 531197
rect 469322 531101 543617 531122
rect 28811 531040 28965 531045
rect 469322 531043 543446 531101
rect 28810 531034 101940 531040
rect 28810 530890 28816 531034
rect 28960 531030 101940 531034
rect 28960 530894 101794 531030
rect 101930 530894 101940 531030
rect 469322 530987 469367 531043
rect 469423 530987 543446 531043
rect 469322 530957 543446 530987
rect 543590 530957 543617 531101
rect 469322 530936 543617 530957
rect 28960 530890 101940 530894
rect 28810 530884 101940 530890
rect 28811 530879 28965 530884
rect 24253 530678 24387 530684
rect 24253 530644 27942 530678
rect 24253 530643 27864 530644
rect 24253 530579 24288 530643
rect 24352 530588 27864 530643
rect 27920 530588 27942 530644
rect 24352 530579 27942 530588
rect 24253 530544 27942 530579
rect 24253 530538 24387 530544
rect -800 507984 19830 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 24593 500484 24711 500490
rect 24593 500457 27734 500484
rect 24593 500393 24620 500457
rect 24684 500452 27734 500457
rect 24684 500396 27660 500452
rect 27716 500396 27734 500452
rect 24684 500393 27734 500396
rect 24593 500366 27734 500393
rect 24593 500360 24711 500366
rect 24913 470292 25031 470298
rect 24913 470265 27734 470292
rect 24913 470201 24940 470265
rect 25004 470260 27734 470265
rect 25004 470204 27660 470260
rect 27716 470204 27734 470260
rect 25004 470201 27734 470204
rect 24913 470174 27734 470201
rect 24913 470168 25031 470174
rect -800 468392 17160 468420
rect -800 468336 17076 468392
rect 17132 468336 17160 468392
rect -800 468308 17160 468336
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 25215 440100 25333 440106
rect 25215 440073 27734 440100
rect 25215 440009 25242 440073
rect 25306 440068 27734 440073
rect 25306 440012 27660 440068
rect 27716 440012 27734 440068
rect 25306 440009 27734 440012
rect 25215 439982 27734 440009
rect 25215 439976 25333 439982
rect -800 425170 22728 425198
rect -800 425114 22644 425170
rect 22700 425114 22728 425170
rect -800 425086 22728 425114
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 25493 409976 25611 409982
rect 25493 409949 27734 409976
rect 25493 409885 25520 409949
rect 25584 409944 27734 409949
rect 25584 409888 27660 409944
rect 27716 409888 27734 409944
rect 25584 409885 27734 409888
rect 25493 409858 27734 409885
rect 25493 409852 25611 409858
rect -800 381948 12344 381976
rect -800 381892 12260 381948
rect 12316 381892 12344 381948
rect -800 381864 12344 381892
rect -800 380682 480 380794
rect 25783 379784 25901 379790
rect 25783 379757 27734 379784
rect 25783 379693 25810 379757
rect 25874 379752 27734 379757
rect 25874 379696 27660 379752
rect 27716 379696 27734 379752
rect 25874 379693 27734 379696
rect 25783 379666 27734 379693
rect 25783 379660 25901 379666
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 26065 349592 26183 349598
rect 26065 349565 27734 349592
rect 26065 349501 26092 349565
rect 26156 349560 27734 349565
rect 26156 349504 27660 349560
rect 27716 349504 27734 349560
rect 26156 349501 27734 349504
rect 26065 349474 27734 349501
rect 26065 349468 26183 349474
rect -800 338726 4710 338754
rect -800 338670 4626 338726
rect 4682 338670 4710 338726
rect -800 338642 4710 338670
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 26317 319468 26435 319474
rect 26317 319441 27734 319468
rect 26317 319377 26344 319441
rect 26408 319436 27734 319441
rect 26408 319380 27660 319436
rect 27716 319380 27734 319436
rect 26408 319377 27734 319380
rect 26317 319350 27734 319377
rect 26317 319344 26435 319350
rect -800 295504 26806 295532
rect -800 295448 26722 295504
rect 26778 295448 26806 295504
rect -800 295420 26806 295448
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect 26554 289666 26674 289700
rect -800 289510 480 289622
rect 26554 289602 26582 289666
rect 26646 289602 26674 289666
rect 26554 289244 26674 289602
rect 26554 289188 26588 289244
rect 26644 289188 26674 289244
rect 26554 289152 26674 289188
rect 544900 269342 547088 582012
rect 550536 313764 552174 587608
rect 552788 530641 553106 530704
rect 552788 530585 552916 530641
rect 552972 530585 553106 530641
rect 552788 530374 553106 530585
rect 552788 530280 552796 530374
rect 552790 530070 552796 530280
rect 553100 530070 553106 530374
rect 552790 530058 553106 530070
rect 556590 358986 558426 611640
rect 563126 405408 563858 617290
rect 568791 449830 569437 621228
rect 573656 494252 574212 623396
rect 577070 583674 577818 627634
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 577070 583562 584800 583674
rect 577070 583558 577818 583562
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 573656 494140 584800 494252
rect 573656 494138 574212 494140
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 568791 449718 584800 449830
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 563126 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 556590 358878 584800 358986
rect 556632 358874 584800 358878
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 550536 313652 584800 313764
rect 583520 275140 584800 275252
rect 555634 274216 555886 274260
rect 555634 274160 555730 274216
rect 555786 274160 555886 274216
rect 555634 273942 555886 274160
rect 583520 273958 584800 274070
rect 555634 273718 555648 273942
rect 555872 273718 555886 273942
rect 555634 273698 555886 273718
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 544900 269230 584800 269342
rect 26784 259263 26914 259302
rect 26784 259199 26817 259263
rect 26881 259199 26914 259263
rect 26784 259052 26914 259199
rect 26784 258996 26820 259052
rect 26876 258996 26914 259052
rect 26784 258976 26914 258996
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248936 14710 248964
rect -800 248880 14626 248936
rect 14682 248880 14710 248936
rect -800 248852 14710 248880
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 27018 229023 27152 229064
rect 27018 228959 27053 229023
rect 27117 228959 27152 229023
rect 27018 228860 27152 228959
rect 27018 228804 27058 228860
rect 27114 228804 27152 228860
rect 27018 228780 27152 228804
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 27246 198945 27380 198986
rect 27246 198881 27281 198945
rect 27345 198881 27380 198945
rect 27246 198736 27380 198881
rect 27246 198680 27286 198736
rect 27342 198680 27380 198736
rect 27246 198662 27380 198680
rect 548619 195130 549289 195135
rect 582340 195130 584800 196230
rect 548618 195106 584800 195130
rect 548618 194482 548642 195106
rect 549266 194482 584800 195106
rect 548618 194458 584800 194482
rect 548619 194453 549289 194458
rect 548673 184250 549343 184255
rect 577294 184250 577966 194458
rect 582340 191430 584800 194458
rect 582340 184250 584800 186230
rect 548672 184226 584800 184250
rect 548672 183602 548696 184226
rect 549320 183602 584800 184226
rect 548672 183578 584800 183602
rect 548673 183573 549343 183578
rect 582340 181430 584800 183578
rect -800 172888 1660 177688
rect 27482 168714 27610 168752
rect 27482 168650 27514 168714
rect 27578 168650 27610 168714
rect 27482 168544 27610 168650
rect 27482 168488 27520 168544
rect 27576 168488 27610 168544
rect 27482 168466 27610 168488
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 27714 138540 27834 138574
rect 27714 138476 27742 138540
rect 27806 138476 27834 138540
rect 27714 138352 27834 138476
rect 27714 138296 27754 138352
rect 27810 138296 27834 138352
rect 27714 138278 27834 138296
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121314 10102 121342
rect -800 121258 10018 121314
rect 10074 121258 10102 121314
rect -800 121230 10102 121258
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 27944 108445 28074 108484
rect 27944 108381 27977 108445
rect 28041 108381 28074 108445
rect 27944 108228 28074 108381
rect 27944 108172 27978 108228
rect 28034 108172 28074 108228
rect 27944 108146 28074 108172
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 580272 92838 584800 92866
rect 580272 92782 580300 92838
rect 580356 92782 584800 92838
rect 580272 92754 584800 92782
rect 583520 91572 584800 91684
rect -800 81638 7272 81666
rect -800 81582 7188 81638
rect 7244 81582 7272 81638
rect -800 81554 7272 81582
rect -800 80372 480 80484
rect -800 79190 480 79302
rect 28176 78506 28340 78522
rect 28176 78362 28186 78506
rect 28330 78362 28340 78506
rect -800 78008 480 78120
rect 28176 78036 28340 78362
rect 28176 77980 28232 78036
rect 28288 77980 28340 78036
rect 28176 77950 28340 77980
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 567598 48180 584800 48208
rect 567598 48124 567626 48180
rect 567682 48124 584800 48180
rect 567598 48096 584800 48124
rect 28482 48065 28640 48078
rect 28482 47921 28489 48065
rect 28633 47921 28640 48065
rect 28482 47844 28640 47921
rect 28482 47788 28524 47844
rect 28580 47788 28640 47844
rect 28482 47752 28640 47788
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect 23608 34898 23720 34904
rect -800 34874 23720 34898
rect -800 34810 23632 34874
rect 23696 34810 23720 34874
rect -800 34786 23720 34810
rect 23608 34780 23720 34786
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 547614 21750 547726 21756
rect 547614 21726 584800 21750
rect 547614 21662 547638 21726
rect 547702 21662 584800 21726
rect 547614 21638 584800 21662
rect 547614 21632 547726 21638
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect 28810 18014 28966 18026
rect 28810 17870 28816 18014
rect 28960 17870 28966 18014
rect 28810 17720 28966 17870
rect 28810 17664 28866 17720
rect 28922 17664 28966 17720
rect 28810 17642 28966 17664
rect 558896 17720 559126 17742
rect 558896 17664 558980 17720
rect 559036 17664 559126 17720
rect 558896 17571 559126 17664
rect 558896 17347 558899 17571
rect 559123 17347 559126 17571
rect 558896 17338 559126 17347
rect 549942 17022 550054 17028
rect -800 16910 480 17022
rect 549942 16998 584800 17022
rect 549942 16934 549966 16998
rect 550030 16934 584800 16998
rect 549942 16910 584800 16934
rect 549942 16904 550054 16910
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect 535055 14918 535725 14923
rect 535054 14894 578558 14918
rect -800 14546 480 14658
rect 535054 14270 535078 14894
rect 535702 14629 578558 14894
rect 535702 14573 578232 14629
rect 578288 14573 578558 14629
rect 535702 14270 578558 14573
rect 582044 14630 584800 14658
rect 582044 14574 582072 14630
rect 582128 14574 584800 14630
rect 582044 14546 584800 14574
rect 535054 14246 578558 14270
rect 535055 14241 535725 14246
rect 22804 13476 22916 13482
rect -800 13452 22916 13476
rect -800 13388 22828 13452
rect 22892 13388 22916 13452
rect -800 13364 22916 13388
rect 22804 13358 22916 13364
rect 552908 13476 553020 13482
rect 552908 13452 584800 13476
rect 552908 13388 552932 13452
rect 552996 13388 584800 13452
rect 552908 13364 584800 13388
rect 552908 13358 553020 13364
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect 582056 9930 583806 9932
rect -800 9818 480 9930
rect 582056 9904 584800 9930
rect 582056 9848 582084 9904
rect 582140 9848 584800 9904
rect 582056 9820 584800 9848
rect 583520 9818 584800 9820
rect 21858 8748 21970 8754
rect -800 8724 21970 8748
rect -800 8660 21882 8724
rect 21946 8660 21970 8724
rect -800 8636 21970 8660
rect 21858 8630 21970 8636
rect 555718 8748 555830 8754
rect 555718 8724 584800 8748
rect 555718 8660 555742 8724
rect 555806 8660 584800 8724
rect 555718 8636 584800 8660
rect 555718 8630 555830 8636
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 582168 5174 584800 5202
rect 582168 5118 582196 5174
rect 582252 5118 584800 5174
rect 582168 5090 584800 5118
rect 20274 4020 20386 4026
rect -800 3996 20386 4020
rect -800 3932 20298 3996
rect 20362 3932 20386 3996
rect -800 3908 20386 3932
rect 20274 3902 20386 3908
rect 558952 4020 559064 4026
rect 558952 3996 584800 4020
rect 558952 3932 558976 3996
rect 559040 3932 584800 3996
rect 558952 3908 584800 3932
rect 558952 3902 559064 3908
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 412672 698801 413216 699345
rect 30438 689933 34822 690797
rect 417408 699226 417712 699235
rect 417408 698931 417412 699226
rect 417412 698931 417708 699226
rect 417708 698931 417712 699226
rect 470570 699226 470874 699235
rect 470570 698931 470574 699226
rect 470574 698931 470870 699226
rect 470870 698931 470874 699226
rect 520606 696782 522990 699166
rect 512854 692664 515238 695048
rect 560058 689678 560362 689687
rect 560058 689383 560062 689678
rect 560062 689383 560358 689678
rect 560358 689383 560362 689678
rect 15022 643920 19646 648544
rect 575946 639838 580650 644542
rect 137844 620284 137988 620428
rect 140294 620284 140438 620428
rect 24288 594466 24352 594530
rect 24620 594172 24684 594236
rect 24940 593876 25004 593940
rect 25242 593608 25306 593672
rect 25520 593338 25584 593402
rect 25810 593026 25874 593090
rect 26092 592736 26156 592800
rect 26344 592446 26408 592510
rect 26582 592176 26646 592240
rect 20222 536797 20446 537021
rect 21680 535600 22144 536064
rect 22694 534572 22998 534876
rect 23520 533513 23824 533817
rect 26817 533082 26881 533146
rect 27053 532840 27117 532904
rect 27281 532590 27345 532654
rect 27514 532346 27578 532410
rect 27742 532128 27806 532192
rect 27977 531868 28041 531932
rect 28186 531536 28330 531680
rect 543448 531365 543592 531509
rect 28489 531204 28633 531348
rect 28816 530890 28960 531034
rect 543446 530957 543590 531101
rect 24288 530579 24352 530643
rect 24620 500393 24684 500457
rect 24940 470201 25004 470265
rect 25242 440009 25306 440073
rect 25520 409885 25584 409949
rect 25810 379693 25874 379757
rect 26092 349501 26156 349565
rect 26344 319377 26408 319441
rect 26582 289602 26646 289666
rect 552796 530070 553100 530374
rect 555648 273718 555872 273942
rect 26817 259199 26881 259263
rect 27053 228959 27117 229023
rect 27281 198881 27345 198945
rect 548642 194482 549266 195106
rect 548696 183602 549320 184226
rect 27514 168650 27578 168714
rect 27742 138476 27806 138540
rect 27977 108381 28041 108445
rect 28186 78362 28330 78506
rect 28489 47921 28633 48065
rect 23632 34810 23696 34874
rect 547638 21662 547702 21726
rect 28816 17870 28960 18014
rect 558899 17347 559123 17571
rect 549966 16934 550030 16998
rect 535078 14270 535702 14894
rect 22828 13388 22892 13452
rect 552932 13388 552996 13452
rect 21882 8660 21946 8724
rect 555742 8660 555806 8724
rect 20298 3932 20362 3996
rect 558976 3932 559040 3996
<< metal4 >>
rect 412640 699376 413248 699377
rect 412640 699345 561426 699376
rect 412640 698801 412672 699345
rect 413216 699235 561426 699345
rect 413216 698931 417408 699235
rect 417712 698931 470570 699235
rect 470874 699204 561426 699235
rect 470874 699166 561436 699204
rect 470874 698931 520606 699166
rect 413216 698801 520606 698931
rect 412640 698770 520606 698801
rect 412640 698769 413248 698770
rect 505280 696782 520606 698770
rect 522990 696782 561436 699166
rect 505280 696744 561436 696782
rect 520567 696743 523029 696744
rect 512815 695048 515277 695087
rect 512815 692664 512854 695048
rect 515238 692664 515277 695048
rect 512815 692625 515277 692664
rect 30276 690797 34940 691006
rect 30276 689933 30438 690797
rect 34822 689933 34940 690797
rect 15001 648564 19667 648565
rect 30276 648564 34940 689933
rect 512816 677318 515276 692625
rect 558976 689687 561436 696744
rect 558976 689383 560058 689687
rect 560362 689383 561436 689687
rect 558976 689304 561436 689383
rect 335440 665430 515346 677318
rect 15001 648544 79422 648564
rect 15001 643920 15022 648544
rect 19646 646916 79422 648544
rect 19646 643920 79482 646916
rect 15001 643900 79482 643920
rect 15001 643899 19667 643900
rect 77850 641872 79482 643900
rect 77850 641072 101504 641872
rect 77850 641066 79482 641072
rect 85622 641066 87254 641072
rect 335440 633052 347328 665430
rect 575937 644550 580659 644551
rect 537992 644546 580659 644550
rect 319632 632252 347328 633052
rect 335440 632248 347328 632252
rect 535732 644542 580659 644546
rect 535732 639838 575946 644542
rect 580650 639838 580659 644542
rect 535732 639830 580659 639838
rect 77850 618834 79482 620798
rect 85622 618834 87254 620798
rect 137840 620431 137992 620432
rect 137840 620428 140441 620431
rect 137840 620284 137844 620428
rect 137988 620284 140294 620428
rect 140438 620284 140441 620428
rect 137840 620281 140441 620284
rect 137840 620280 137992 620281
rect 24253 594530 24387 594565
rect 24253 594466 24288 594530
rect 24352 594466 24387 594530
rect 20194 537021 20474 537049
rect 20194 536797 20222 537021
rect 20446 536797 20474 537021
rect 20194 536769 20474 536797
rect 20195 3996 20473 536769
rect 21651 536064 22173 536093
rect 21651 535600 21680 536064
rect 22144 535600 22173 536064
rect 21651 535571 22173 535600
rect 21652 8724 22172 535571
rect 22675 534876 23017 534895
rect 22675 534572 22694 534876
rect 22998 534572 23017 534876
rect 22675 534553 23017 534572
rect 22676 13452 23016 534553
rect 23488 533817 23856 533849
rect 23488 533513 23520 533817
rect 23824 533513 23856 533817
rect 23488 533481 23856 533513
rect 23489 34874 23855 533481
rect 24253 530679 24387 594466
rect 24593 594236 24711 594263
rect 24593 594172 24620 594236
rect 24684 594172 24711 594236
rect 24252 530643 24388 530679
rect 24252 530579 24288 530643
rect 24352 530579 24388 530643
rect 24252 530543 24388 530579
rect 24593 500485 24711 594172
rect 24913 593940 25031 593967
rect 24913 593876 24940 593940
rect 25004 593876 25031 593940
rect 24592 500457 24712 500485
rect 24592 500393 24620 500457
rect 24684 500393 24712 500457
rect 24592 500365 24712 500393
rect 24913 470293 25031 593876
rect 25215 593672 25333 593699
rect 25215 593608 25242 593672
rect 25306 593608 25333 593672
rect 24912 470265 25032 470293
rect 24912 470201 24940 470265
rect 25004 470201 25032 470265
rect 24912 470173 25032 470201
rect 25215 440101 25333 593608
rect 25493 593402 25611 593429
rect 25493 593338 25520 593402
rect 25584 593338 25611 593402
rect 25214 440073 25334 440101
rect 25214 440009 25242 440073
rect 25306 440009 25334 440073
rect 25214 439981 25334 440009
rect 25493 409977 25611 593338
rect 25783 593090 25901 593117
rect 25783 593026 25810 593090
rect 25874 593026 25901 593090
rect 25492 409949 25612 409977
rect 25492 409885 25520 409949
rect 25584 409885 25612 409949
rect 25492 409857 25612 409885
rect 25783 379785 25901 593026
rect 26065 592800 26183 592827
rect 26065 592736 26092 592800
rect 26156 592736 26183 592800
rect 25782 379757 25902 379785
rect 25782 379693 25810 379757
rect 25874 379693 25902 379757
rect 25782 379665 25902 379693
rect 26065 349593 26183 592736
rect 26317 592510 26435 592537
rect 26317 592446 26344 592510
rect 26408 592446 26435 592510
rect 26064 349565 26184 349593
rect 26064 349501 26092 349565
rect 26156 349501 26184 349565
rect 26064 349473 26184 349501
rect 26317 319469 26435 592446
rect 26554 592240 26674 592268
rect 26554 592176 26582 592240
rect 26646 592176 26674 592240
rect 26316 319441 26436 319469
rect 26316 319377 26344 319441
rect 26408 319377 26436 319441
rect 26316 319349 26436 319377
rect 26554 289695 26674 592176
rect 75402 566818 77034 607942
rect 77850 600360 79482 605350
rect 85622 600360 87254 605302
rect 77848 599560 87254 600360
rect 77850 567218 79482 599560
rect 85622 568074 87254 599560
rect 88070 568472 89702 607942
rect 75418 534000 77050 556592
rect 77866 549010 79498 554000
rect 85638 549010 87270 553952
rect 77864 548210 87270 549010
rect 26784 533146 26914 533179
rect 26784 533082 26817 533146
rect 26881 533082 26914 533146
rect 26553 289666 26675 289695
rect 26553 289602 26582 289666
rect 26646 289602 26675 289666
rect 26553 289573 26675 289602
rect 26784 259297 26914 533082
rect 27018 532904 27152 532939
rect 27018 532840 27053 532904
rect 27117 532840 27152 532904
rect 26783 259263 26915 259297
rect 26783 259199 26817 259263
rect 26881 259199 26915 259263
rect 26783 259165 26915 259199
rect 27018 229059 27152 532840
rect 27246 532654 27380 532689
rect 27246 532590 27281 532654
rect 27345 532590 27380 532654
rect 27017 229023 27153 229059
rect 27017 228959 27053 229023
rect 27117 228959 27153 229023
rect 27017 228923 27153 228959
rect 27246 198981 27380 532590
rect 27482 532410 27610 532442
rect 27482 532346 27514 532410
rect 27578 532346 27610 532410
rect 75418 532368 78776 534000
rect 27245 198945 27381 198981
rect 27245 198881 27281 198945
rect 27345 198881 27381 198945
rect 27245 198845 27381 198881
rect 27482 168747 27610 532346
rect 27714 532192 27834 532220
rect 27714 532128 27742 532192
rect 27806 532128 27834 532192
rect 27481 168714 27611 168747
rect 27481 168650 27514 168714
rect 27578 168650 27611 168714
rect 27481 168617 27611 168650
rect 27714 138569 27834 532128
rect 27944 531932 28074 531965
rect 27944 531868 27977 531932
rect 28041 531868 28074 531932
rect 27713 138540 27835 138569
rect 27713 138476 27742 138540
rect 27806 138476 27835 138540
rect 27713 138447 27835 138476
rect 27944 108479 28074 531868
rect 28176 531680 28340 531690
rect 28176 531536 28186 531680
rect 28330 531536 28340 531680
rect 27943 108445 28075 108479
rect 27943 108381 27977 108445
rect 28041 108381 28075 108445
rect 27943 108347 28075 108381
rect 28176 78517 28340 531536
rect 28482 531348 28640 531355
rect 28482 531204 28489 531348
rect 28633 531204 28640 531348
rect 28175 78506 28341 78517
rect 28175 78362 28186 78506
rect 28330 78362 28341 78506
rect 28175 78351 28341 78362
rect 28482 48073 28640 531204
rect 28810 531034 28966 531040
rect 28810 530890 28816 531034
rect 28960 530890 28966 531034
rect 28481 48065 28641 48073
rect 28481 47921 28489 48065
rect 28633 47921 28641 48065
rect 28481 47913 28641 47921
rect 23489 34810 23632 34874
rect 23696 34810 23855 34874
rect 23489 34720 23855 34810
rect 28810 18021 28966 530890
rect 78094 500366 78766 532368
rect 80746 531852 81546 548210
rect 88086 532276 89718 554700
rect 535732 532446 541064 639830
rect 575937 639829 580659 639830
rect 80814 496902 81486 531852
rect 88974 504554 89646 532276
rect 537882 510238 539514 532446
rect 543418 531538 543622 531539
rect 543418 531509 550107 531538
rect 543418 531365 543448 531509
rect 543592 531365 550107 531509
rect 543418 531336 550107 531365
rect 543418 531335 543622 531336
rect 543424 531122 543612 531123
rect 543424 531101 547764 531122
rect 543424 530957 543446 531101
rect 543590 530957 547764 531101
rect 543424 530936 547764 530957
rect 543424 530935 543612 530936
rect 28809 18014 28967 18021
rect 28809 17870 28816 18014
rect 28960 17870 28967 18014
rect 28809 17863 28967 17870
rect 535054 14894 535726 39862
rect 547578 21726 547764 530936
rect 548618 195106 549290 195130
rect 548618 194482 548642 195106
rect 549266 194482 549290 195106
rect 548618 194458 549290 194482
rect 548672 184226 549344 184250
rect 548672 183602 548696 184226
rect 549320 183602 549344 184226
rect 548672 183578 549344 183602
rect 547578 21662 547638 21726
rect 547702 21662 547764 21726
rect 547578 21599 547764 21662
rect 549905 16998 550107 531336
rect 552789 530380 553107 530381
rect 549905 16934 549966 16998
rect 550030 16934 550107 16998
rect 549905 16879 550107 16934
rect 552784 530374 553110 530380
rect 552784 530070 552796 530374
rect 553100 530206 553110 530374
rect 553100 530070 553112 530206
rect 535054 14270 535078 14894
rect 535702 14270 535726 14894
rect 535054 14246 535726 14270
rect 22676 13388 22828 13452
rect 22892 13388 23016 13452
rect 22676 13346 23016 13388
rect 552784 13452 553112 530070
rect 555633 273942 555887 273957
rect 555633 273718 555648 273942
rect 555872 273718 555887 273942
rect 555633 273703 555887 273718
rect 552784 13388 552932 13452
rect 552996 13388 553112 13452
rect 552784 13322 553112 13388
rect 21652 8660 21882 8724
rect 21946 8660 22172 8724
rect 21652 8596 22172 8660
rect 555634 8724 555886 273703
rect 558895 17571 559127 17575
rect 558895 17347 558899 17571
rect 559123 17347 559127 17571
rect 558895 17343 559127 17347
rect 555634 8660 555742 8724
rect 555806 8660 555886 8724
rect 555634 8596 555886 8660
rect 20195 3932 20298 3996
rect 20362 3932 20473 3996
rect 20195 3871 20473 3932
rect 558896 3996 559126 17343
rect 558896 3932 558976 3996
rect 559040 3932 559126 3996
rect 558896 3869 559126 3932
<< via4 >>
rect 548676 194516 549232 195072
rect 548730 183636 549286 184192
<< metal5 >>
rect 93520 621340 93548 621350
rect 539778 195072 549290 195130
rect 539778 194516 548676 195072
rect 549232 194516 549290 195072
rect 539778 194458 549290 194516
rect 540754 184192 549344 184250
rect 540754 183636 548730 184192
rect 549286 183636 549344 184192
rect 540754 183578 549344 183636
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_6
timestamp 1624302123
transform 0 1 579599 -1 0 14602
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_7
timestamp 1624302123
transform 0 1 579611 -1 0 9876
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_8
timestamp 1624302123
transform 0 1 579723 -1 0 5146
box -60 -357 60 357
use analog_top_level  analog_top_level_0
timestamp 1624302123
transform -1 0 479200 0 1 739592
box 157324 -188462 385680 -59028
use sar_adc_controller_8bit  sar_adc_controller_8bit_1
timestamp 1624302123
transform -1 0 90618 0 -1 570806
box 0 0 16100 20128
use sar_adc_controller_8bit  sar_adc_controller_8bit_0
timestamp 1624302123
transform -1 0 90602 0 -1 622156
box 0 0 16100 20128
use esd_cell  esd_cell_10
timestamp 1624302123
transform 1 0 5996 0 1 682782
box -2400 -3178 2400 3178
use esd_cell  esd_cell_9
timestamp 1624302123
transform 1 0 22248 0 1 697476
box -2400 -3178 2400 3178
use esd_cell  esd_cell_8
timestamp 1624302123
transform 1 0 75404 0 1 697476
box -2400 -3178 2400 3178
use esd_cell  esd_cell_7
timestamp 1624302123
transform 1 0 127332 0 1 698616
box -2400 -3178 2400 3178
use esd_cell  esd_cell_6
timestamp 1624302123
transform 1 0 215186 0 1 695212
box -2400 -3178 2400 3178
use esd_cell  esd_cell_5
timestamp 1624302123
transform 1 0 200032 0 1 689638
box -2400 -3178 2400 3178
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_4
timestamp 1624302123
transform -1 0 171964 0 -1 701565
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_5
timestamp 1624302123
transform -1 0 174470 0 -1 701565
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_2
timestamp 1624302123
transform -1 0 226152 0 -1 701565
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_3
timestamp 1624302123
transform -1 0 223752 0 -1 701565
box -60 -357 60 357
use esd_cell  esd_cell_4
timestamp 1624302123
transform 1 0 408838 0 1 696756
box -2400 -3178 2400 3178
use esd_cell  esd_cell_3
timestamp 1624302123
transform 1 0 318206 0 1 694824
box -2400 -3178 2400 3178
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_1
timestamp 1624302123
transform -1 0 327900 0 -1 701565
box -60 -357 60 357
use sky130_fd_pr__res_generic_m1_DYSWBR  sky130_fd_pr__res_generic_m1_DYSWBR_0
timestamp 1624302123
transform -1 0 325390 0 -1 701565
box -60 -357 60 357
use esd_cell  esd_cell_2
timestamp 1624302123
transform 1 0 463684 0 1 693044
box -2400 -3178 2400 3178
use esd_cell  esd_cell_1
timestamp 1624302123
transform 1 0 577108 0 1 680432
box -2400 -3178 2400 3178
use esd_cell  esd_cell_0
timestamp 1624302123
transform 1 0 566444 0 1 692528
box -2400 -3178 2400 3178
use deconv_kernel_estimator_top_level  deconv_kernel_estimator_top_level_0
timestamp 1624302123
transform 1 0 29134 0 1 17658
box 0 0 513728 512992
<< labels >>
flabel metal3 s 97138 619918 97180 619954 1 FreeSans 600 0 0 0 sig_frequency_7
flabel metal3 s 97036 617672 97078 617714 1 FreeSans 600 0 0 0 sig_frequency_6
flabel metal3 s 96998 615414 97028 615456 1 FreeSans 600 0 0 0 sig_frequency_5
flabel metal3 s 96882 613170 96918 613214 1 FreeSans 600 0 0 0 sig_frequency_4
flabel metal3 s 96900 610990 96924 611028 1 FreeSans 600 0 0 0 sig_frequency_3
flabel metal3 s 96764 608770 96790 608796 1 FreeSans 600 0 0 0 sig_frequency_2
flabel metal3 s 96722 606516 96752 606564 1 FreeSans 600 0 0 0 sig_frequency_1
flabel metal3 s 96746 604278 96802 604328 1 FreeSans 600 0 0 0 sig_frequency_0
flabel metal3 s 137200 620356 137222 620376 1 FreeSans 600 0 0 0 sample
flabel metal3 s 97254 552942 97336 552992 1 FreeSans 600 0 0 0 sig_amplitude_0
flabel metal3 s 97126 555166 97172 555212 1 FreeSans 600 0 0 0 sig_amplitude_1
flabel metal3 s 96984 557436 97020 557470 1 FreeSans 600 0 0 0 sig_amplitude_2
flabel metal3 s 96762 559642 96798 559674 1 FreeSans 600 0 0 0 sig_amplitude_3
flabel metal3 s 96656 561850 96696 561878 1 FreeSans 600 0 0 0 sig_amplitude_4
flabel metal3 s 96516 564072 96548 564108 1 FreeSans 600 0 0 0 sig_amplitude_5
flabel metal3 s 96390 566330 96434 566374 1 FreeSans 600 0 0 0 sig_amplitude_6
flabel metal3 s 96328 567996 96364 568042 1 FreeSans 600 0 0 0 sig_amplitude_7
flabel metal2 s 92812 587564 92830 587588 1 FreeSans 600 0 0 0 amplitude_comparator_val
flabel metal2 s 92824 638576 92846 638598 1 FreeSans 600 0 0 0 frequency_comparator_val
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1750 0 0 0 gpio_analog[0]
port 1 nsew
flabel metal3 s -800 381864 480 381976 0 FreeSans 1750 0 0 0 gpio_analog[10]
port 2 nsew
flabel metal3 s -800 338642 480 338754 0 FreeSans 1750 0 0 0 gpio_analog[11]
port 3 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1750 0 0 0 gpio_analog[12]
port 4 nsew
flabel metal3 s -800 252398 480 252510 0 FreeSans 1750 0 0 0 gpio_analog[13]
port 5 nsew
flabel metal3 s -800 124776 480 124888 0 FreeSans 1750 0 0 0 gpio_analog[14]
port 6 nsew
flabel metal3 s -800 81554 480 81666 0 FreeSans 1750 0 0 0 gpio_analog[15]
port 7 nsew
flabel metal3 s -800 38332 480 38444 0 FreeSans 1750 0 0 0 gpio_analog[16]
port 8 nsew
flabel metal3 s -800 16910 480 17022 0 FreeSans 1750 0 0 0 gpio_analog[17]
port 9 nsew
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1750 0 0 0 gpio_analog[1]
port 10 nsew
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1750 0 0 0 gpio_analog[2]
port 11 nsew
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1750 0 0 0 gpio_analog[3]
port 12 nsew
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1750 0 0 0 gpio_analog[4]
port 13 nsew
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1750 0 0 0 gpio_analog[5]
port 14 nsew
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1750 0 0 0 gpio_analog[6]
port 15 nsew
flabel metal3 s -800 511530 480 511642 0 FreeSans 1750 0 0 0 gpio_analog[7]
port 16 nsew
flabel metal3 s -800 468308 480 468420 0 FreeSans 1750 0 0 0 gpio_analog[8]
port 17 nsew
flabel metal3 s -800 425086 480 425198 0 FreeSans 1750 0 0 0 gpio_analog[9]
port 18 nsew
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1750 0 0 0 gpio_noesd[0]
port 19 nsew
flabel metal3 s -800 380682 480 380794 0 FreeSans 1750 0 0 0 gpio_noesd[10]
port 20 nsew
flabel metal3 s -800 337460 480 337572 0 FreeSans 1750 0 0 0 gpio_noesd[11]
port 21 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1750 0 0 0 gpio_noesd[12]
port 22 nsew
flabel metal3 s -800 251216 480 251328 0 FreeSans 1750 0 0 0 gpio_noesd[13]
port 23 nsew
flabel metal3 s -800 123594 480 123706 0 FreeSans 1750 0 0 0 gpio_noesd[14]
port 24 nsew
flabel metal3 s -800 80372 480 80484 0 FreeSans 1750 0 0 0 gpio_noesd[15]
port 25 nsew
flabel metal3 s -800 37150 480 37262 0 FreeSans 1750 0 0 0 gpio_noesd[16]
port 26 nsew
flabel metal3 s -800 15728 480 15840 0 FreeSans 1750 0 0 0 gpio_noesd[17]
port 27 nsew
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1750 0 0 0 gpio_noesd[1]
port 28 nsew
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1750 0 0 0 gpio_noesd[2]
port 29 nsew
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1750 0 0 0 gpio_noesd[3]
port 30 nsew
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1750 0 0 0 gpio_noesd[4]
port 31 nsew
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1750 0 0 0 gpio_noesd[5]
port 32 nsew
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1750 0 0 0 gpio_noesd[6]
port 33 nsew
flabel metal3 s -800 510348 480 510460 0 FreeSans 1750 0 0 0 gpio_noesd[7]
port 34 nsew
flabel metal3 s -800 467126 480 467238 0 FreeSans 1750 0 0 0 gpio_noesd[8]
port 35 nsew
flabel metal3 s -800 423904 480 424016 0 FreeSans 1750 0 0 0 gpio_noesd[9]
port 36 nsew
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1750 0 0 0 io_analog[0]
port 37 nsew
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1750 0 0 0 io_analog[10]
port 38 nsew
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 3000 180 0 0 io_analog[1]
port 39 nsew
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 3000 180 0 0 io_analog[2]
port 40 nsew
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 3000 180 0 0 io_analog[3]
port 41 nsew
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 3000 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 3000 180 0 0 io_analog[4]
port 42 nsew
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 3000 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 3000 180 0 0 io_analog[5]
port 43 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 3000 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 3000 180 0 0 io_analog[6]
port 44 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 3000 180 0 0 io_analog[7]
port 45 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 3000 180 0 0 io_analog[8]
port 46 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 3000 180 0 0 io_analog[9]
port 47 nsew
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 3000 180 0 0 io_clamp_high[0]
port 48 nsew
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 3000 180 0 0 io_clamp_high[1]
port 49 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 3000 180 0 0 io_clamp_high[2]
port 50 nsew
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 3000 180 0 0 io_clamp_low[0]
port 51 nsew
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 3000 180 0 0 io_clamp_low[1]
port 52 nsew
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 3000 180 0 0 io_clamp_low[2]
port 53 nsew
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1750 0 0 0 io_in[0]
port 54 nsew
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1750 0 0 0 io_in[10]
port 55 nsew
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1750 0 0 0 io_in[11]
port 56 nsew
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1750 0 0 0 io_in[12]
port 57 nsew
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1750 0 0 0 io_in[13]
port 58 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1750 0 0 0 io_in[14]
port 59 nsew
flabel metal3 s -800 464762 480 464874 0 FreeSans 1750 0 0 0 io_in[15]
port 60 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1750 0 0 0 io_in[16]
port 61 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1750 0 0 0 io_in[17]
port 62 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1750 0 0 0 io_in[18]
port 63 nsew
flabel metal3 s -800 291874 480 291986 0 FreeSans 1750 0 0 0 io_in[19]
port 64 nsew
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1750 0 0 0 io_in[1]
port 65 nsew
flabel metal3 s -800 248852 480 248964 0 FreeSans 1750 0 0 0 io_in[20]
port 66 nsew
flabel metal3 s -800 121230 480 121342 0 FreeSans 1750 0 0 0 io_in[21]
port 67 nsew
flabel metal3 s -800 78008 480 78120 0 FreeSans 1750 0 0 0 io_in[22]
port 68 nsew
flabel metal3 s -800 34786 480 34898 0 FreeSans 1750 0 0 0 io_in[23]
port 69 nsew
flabel metal3 s -800 13364 480 13476 0 FreeSans 1750 0 0 0 io_in[24]
port 70 nsew
flabel metal3 s -800 8636 480 8748 0 FreeSans 1750 0 0 0 io_in[25]
port 71 nsew
flabel metal3 s -800 3908 480 4020 0 FreeSans 1750 0 0 0 io_in[26]
port 72 nsew
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1750 0 0 0 io_in[2]
port 73 nsew
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1750 0 0 0 io_in[3]
port 74 nsew
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1750 0 0 0 io_in[4]
port 75 nsew
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1750 0 0 0 io_in[5]
port 76 nsew
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1750 0 0 0 io_in[6]
port 77 nsew
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1750 0 0 0 io_in[7]
port 78 nsew
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1750 0 0 0 io_in[8]
port 79 nsew
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1750 0 0 0 io_in[9]
port 80 nsew
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1750 0 0 0 io_in_3v3[0]
port 81 nsew
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1750 0 0 0 io_in_3v3[10]
port 82 nsew
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1750 0 0 0 io_in_3v3[11]
port 83 nsew
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1750 0 0 0 io_in_3v3[12]
port 84 nsew
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1750 0 0 0 io_in_3v3[13]
port 85 nsew
flabel metal3 s -800 509166 480 509278 0 FreeSans 1750 0 0 0 io_in_3v3[14]
port 86 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1750 0 0 0 io_in_3v3[15]
port 87 nsew
flabel metal3 s -800 422722 480 422834 0 FreeSans 1750 0 0 0 io_in_3v3[16]
port 88 nsew
flabel metal3 s -800 379500 480 379612 0 FreeSans 1750 0 0 0 io_in_3v3[17]
port 89 nsew
flabel metal3 s -800 336278 480 336390 0 FreeSans 1750 0 0 0 io_in_3v3[18]
port 90 nsew
flabel metal3 s -800 293056 480 293168 0 FreeSans 1750 0 0 0 io_in_3v3[19]
port 91 nsew
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1750 0 0 0 io_in_3v3[1]
port 92 nsew
flabel metal3 s -800 250034 480 250146 0 FreeSans 1750 0 0 0 io_in_3v3[20]
port 93 nsew
flabel metal3 s -800 122412 480 122524 0 FreeSans 1750 0 0 0 io_in_3v3[21]
port 94 nsew
flabel metal3 s -800 79190 480 79302 0 FreeSans 1750 0 0 0 io_in_3v3[22]
port 95 nsew
flabel metal3 s -800 35968 480 36080 0 FreeSans 1750 0 0 0 io_in_3v3[23]
port 96 nsew
flabel metal3 s -800 14546 480 14658 0 FreeSans 1750 0 0 0 io_in_3v3[24]
port 97 nsew
flabel metal3 s -800 9818 480 9930 0 FreeSans 1750 0 0 0 io_in_3v3[25]
port 98 nsew
flabel metal3 s -800 5090 480 5202 0 FreeSans 1750 0 0 0 io_in_3v3[26]
port 99 nsew
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1750 0 0 0 io_in_3v3[2]
port 100 nsew
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1750 0 0 0 io_in_3v3[3]
port 101 nsew
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1750 0 0 0 io_in_3v3[4]
port 102 nsew
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1750 0 0 0 io_in_3v3[5]
port 103 nsew
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1750 0 0 0 io_in_3v3[6]
port 104 nsew
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1750 0 0 0 io_in_3v3[7]
port 105 nsew
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1750 0 0 0 io_in_3v3[8]
port 106 nsew
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1750 0 0 0 io_in_3v3[9]
port 107 nsew
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1750 0 0 0 io_oeb[0]
port 108 nsew
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1750 0 0 0 io_oeb[10]
port 109 nsew
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1750 0 0 0 io_oeb[11]
port 110 nsew
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1750 0 0 0 io_oeb[12]
port 111 nsew
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1750 0 0 0 io_oeb[13]
port 112 nsew
flabel metal3 s -800 505620 480 505732 0 FreeSans 1750 0 0 0 io_oeb[14]
port 113 nsew
flabel metal3 s -800 462398 480 462510 0 FreeSans 1750 0 0 0 io_oeb[15]
port 114 nsew
flabel metal3 s -800 419176 480 419288 0 FreeSans 1750 0 0 0 io_oeb[16]
port 115 nsew
flabel metal3 s -800 375954 480 376066 0 FreeSans 1750 0 0 0 io_oeb[17]
port 116 nsew
flabel metal3 s -800 332732 480 332844 0 FreeSans 1750 0 0 0 io_oeb[18]
port 117 nsew
flabel metal3 s -800 289510 480 289622 0 FreeSans 1750 0 0 0 io_oeb[19]
port 118 nsew
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1750 0 0 0 io_oeb[1]
port 119 nsew
flabel metal3 s -800 246488 480 246600 0 FreeSans 1750 0 0 0 io_oeb[20]
port 120 nsew
flabel metal3 s -800 118866 480 118978 0 FreeSans 1750 0 0 0 io_oeb[21]
port 121 nsew
flabel metal3 s -800 75644 480 75756 0 FreeSans 1750 0 0 0 io_oeb[22]
port 122 nsew
flabel metal3 s -800 32422 480 32534 0 FreeSans 1750 0 0 0 io_oeb[23]
port 123 nsew
flabel metal3 s -800 11000 480 11112 0 FreeSans 1750 0 0 0 io_oeb[24]
port 124 nsew
flabel metal3 s -800 6272 480 6384 0 FreeSans 1750 0 0 0 io_oeb[25]
port 125 nsew
flabel metal3 s -800 1544 480 1656 0 FreeSans 1750 0 0 0 io_oeb[26]
port 126 nsew
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1750 0 0 0 io_oeb[2]
port 127 nsew
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1750 0 0 0 io_oeb[3]
port 128 nsew
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1750 0 0 0 io_oeb[4]
port 129 nsew
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1750 0 0 0 io_oeb[5]
port 130 nsew
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1750 0 0 0 io_oeb[6]
port 131 nsew
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1750 0 0 0 io_oeb[7]
port 132 nsew
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1750 0 0 0 io_oeb[8]
port 133 nsew
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1750 0 0 0 io_oeb[9]
port 134 nsew
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1750 0 0 0 io_out[0]
port 135 nsew
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1750 0 0 0 io_out[10]
port 136 nsew
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1750 0 0 0 io_out[11]
port 137 nsew
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1750 0 0 0 io_out[12]
port 138 nsew
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1750 0 0 0 io_out[13]
port 139 nsew
flabel metal3 s -800 506802 480 506914 0 FreeSans 1750 0 0 0 io_out[14]
port 140 nsew
flabel metal3 s -800 463580 480 463692 0 FreeSans 1750 0 0 0 io_out[15]
port 141 nsew
flabel metal3 s -800 420358 480 420470 0 FreeSans 1750 0 0 0 io_out[16]
port 142 nsew
flabel metal3 s -800 377136 480 377248 0 FreeSans 1750 0 0 0 io_out[17]
port 143 nsew
flabel metal3 s -800 333914 480 334026 0 FreeSans 1750 0 0 0 io_out[18]
port 144 nsew
flabel metal3 s -800 290692 480 290804 0 FreeSans 1750 0 0 0 io_out[19]
port 145 nsew
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1750 0 0 0 io_out[1]
port 146 nsew
flabel metal3 s -800 247670 480 247782 0 FreeSans 1750 0 0 0 io_out[20]
port 147 nsew
flabel metal3 s -800 120048 480 120160 0 FreeSans 1750 0 0 0 io_out[21]
port 148 nsew
flabel metal3 s -800 76826 480 76938 0 FreeSans 1750 0 0 0 io_out[22]
port 149 nsew
flabel metal3 s -800 33604 480 33716 0 FreeSans 1750 0 0 0 io_out[23]
port 150 nsew
flabel metal3 s -800 12182 480 12294 0 FreeSans 1750 0 0 0 io_out[24]
port 151 nsew
flabel metal3 s -800 7454 480 7566 0 FreeSans 1750 0 0 0 io_out[25]
port 152 nsew
flabel metal3 s -800 2726 480 2838 0 FreeSans 1750 0 0 0 io_out[26]
port 153 nsew
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1750 0 0 0 io_out[2]
port 154 nsew
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1750 0 0 0 io_out[3]
port 155 nsew
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1750 0 0 0 io_out[4]
port 156 nsew
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1750 0 0 0 io_out[5]
port 157 nsew
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1750 0 0 0 io_out[6]
port 158 nsew
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1750 0 0 0 io_out[7]
port 159 nsew
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1750 0 0 0 io_out[8]
port 160 nsew
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1750 0 0 0 io_out[9]
port 161 nsew
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1750 90 0 0 la_data_in[0]
port 162 nsew
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1750 90 0 0 la_data_in[100]
port 163 nsew
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1750 90 0 0 la_data_in[101]
port 164 nsew
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1750 90 0 0 la_data_in[102]
port 165 nsew
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1750 90 0 0 la_data_in[103]
port 166 nsew
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1750 90 0 0 la_data_in[104]
port 167 nsew
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1750 90 0 0 la_data_in[105]
port 168 nsew
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1750 90 0 0 la_data_in[106]
port 169 nsew
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1750 90 0 0 la_data_in[107]
port 170 nsew
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1750 90 0 0 la_data_in[108]
port 171 nsew
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1750 90 0 0 la_data_in[109]
port 172 nsew
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1750 90 0 0 la_data_in[10]
port 173 nsew
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1750 90 0 0 la_data_in[110]
port 174 nsew
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1750 90 0 0 la_data_in[111]
port 175 nsew
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1750 90 0 0 la_data_in[112]
port 176 nsew
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1750 90 0 0 la_data_in[113]
port 177 nsew
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1750 90 0 0 la_data_in[114]
port 178 nsew
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1750 90 0 0 la_data_in[115]
port 179 nsew
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1750 90 0 0 la_data_in[116]
port 180 nsew
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1750 90 0 0 la_data_in[117]
port 181 nsew
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1750 90 0 0 la_data_in[118]
port 182 nsew
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1750 90 0 0 la_data_in[119]
port 183 nsew
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1750 90 0 0 la_data_in[11]
port 184 nsew
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1750 90 0 0 la_data_in[120]
port 185 nsew
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1750 90 0 0 la_data_in[121]
port 186 nsew
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1750 90 0 0 la_data_in[122]
port 187 nsew
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1750 90 0 0 la_data_in[123]
port 188 nsew
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1750 90 0 0 la_data_in[124]
port 189 nsew
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1750 90 0 0 la_data_in[125]
port 190 nsew
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1750 90 0 0 la_data_in[126]
port 191 nsew
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1750 90 0 0 la_data_in[127]
port 192 nsew
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1750 90 0 0 la_data_in[12]
port 193 nsew
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1750 90 0 0 la_data_in[13]
port 194 nsew
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1750 90 0 0 la_data_in[14]
port 195 nsew
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1750 90 0 0 la_data_in[15]
port 196 nsew
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1750 90 0 0 la_data_in[16]
port 197 nsew
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1750 90 0 0 la_data_in[17]
port 198 nsew
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1750 90 0 0 la_data_in[18]
port 199 nsew
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1750 90 0 0 la_data_in[19]
port 200 nsew
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1750 90 0 0 la_data_in[1]
port 201 nsew
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1750 90 0 0 la_data_in[20]
port 202 nsew
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1750 90 0 0 la_data_in[21]
port 203 nsew
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1750 90 0 0 la_data_in[22]
port 204 nsew
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1750 90 0 0 la_data_in[23]
port 205 nsew
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1750 90 0 0 la_data_in[24]
port 206 nsew
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1750 90 0 0 la_data_in[25]
port 207 nsew
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1750 90 0 0 la_data_in[26]
port 208 nsew
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1750 90 0 0 la_data_in[27]
port 209 nsew
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1750 90 0 0 la_data_in[28]
port 210 nsew
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1750 90 0 0 la_data_in[29]
port 211 nsew
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1750 90 0 0 la_data_in[2]
port 212 nsew
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1750 90 0 0 la_data_in[30]
port 213 nsew
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1750 90 0 0 la_data_in[31]
port 214 nsew
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1750 90 0 0 la_data_in[32]
port 215 nsew
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1750 90 0 0 la_data_in[33]
port 216 nsew
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1750 90 0 0 la_data_in[34]
port 217 nsew
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1750 90 0 0 la_data_in[35]
port 218 nsew
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1750 90 0 0 la_data_in[36]
port 219 nsew
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1750 90 0 0 la_data_in[37]
port 220 nsew
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1750 90 0 0 la_data_in[38]
port 221 nsew
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1750 90 0 0 la_data_in[39]
port 222 nsew
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1750 90 0 0 la_data_in[3]
port 223 nsew
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1750 90 0 0 la_data_in[40]
port 224 nsew
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1750 90 0 0 la_data_in[41]
port 225 nsew
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1750 90 0 0 la_data_in[42]
port 226 nsew
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1750 90 0 0 la_data_in[43]
port 227 nsew
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1750 90 0 0 la_data_in[44]
port 228 nsew
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1750 90 0 0 la_data_in[45]
port 229 nsew
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1750 90 0 0 la_data_in[46]
port 230 nsew
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1750 90 0 0 la_data_in[47]
port 231 nsew
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1750 90 0 0 la_data_in[48]
port 232 nsew
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1750 90 0 0 la_data_in[49]
port 233 nsew
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1750 90 0 0 la_data_in[4]
port 234 nsew
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1750 90 0 0 la_data_in[50]
port 235 nsew
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1750 90 0 0 la_data_in[51]
port 236 nsew
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1750 90 0 0 la_data_in[52]
port 237 nsew
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1750 90 0 0 la_data_in[53]
port 238 nsew
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1750 90 0 0 la_data_in[54]
port 239 nsew
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1750 90 0 0 la_data_in[55]
port 240 nsew
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1750 90 0 0 la_data_in[56]
port 241 nsew
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1750 90 0 0 la_data_in[57]
port 242 nsew
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1750 90 0 0 la_data_in[58]
port 243 nsew
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1750 90 0 0 la_data_in[59]
port 244 nsew
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1750 90 0 0 la_data_in[5]
port 245 nsew
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1750 90 0 0 la_data_in[60]
port 246 nsew
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1750 90 0 0 la_data_in[61]
port 247 nsew
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1750 90 0 0 la_data_in[62]
port 248 nsew
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1750 90 0 0 la_data_in[63]
port 249 nsew
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1750 90 0 0 la_data_in[64]
port 250 nsew
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1750 90 0 0 la_data_in[65]
port 251 nsew
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1750 90 0 0 la_data_in[66]
port 252 nsew
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1750 90 0 0 la_data_in[67]
port 253 nsew
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1750 90 0 0 la_data_in[68]
port 254 nsew
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1750 90 0 0 la_data_in[69]
port 255 nsew
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1750 90 0 0 la_data_in[6]
port 256 nsew
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1750 90 0 0 la_data_in[70]
port 257 nsew
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1750 90 0 0 la_data_in[71]
port 258 nsew
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1750 90 0 0 la_data_in[72]
port 259 nsew
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1750 90 0 0 la_data_in[73]
port 260 nsew
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1750 90 0 0 la_data_in[74]
port 261 nsew
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1750 90 0 0 la_data_in[75]
port 262 nsew
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1750 90 0 0 la_data_in[76]
port 263 nsew
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1750 90 0 0 la_data_in[77]
port 264 nsew
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1750 90 0 0 la_data_in[78]
port 265 nsew
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1750 90 0 0 la_data_in[79]
port 266 nsew
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1750 90 0 0 la_data_in[7]
port 267 nsew
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1750 90 0 0 la_data_in[80]
port 268 nsew
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1750 90 0 0 la_data_in[81]
port 269 nsew
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1750 90 0 0 la_data_in[82]
port 270 nsew
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1750 90 0 0 la_data_in[83]
port 271 nsew
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1750 90 0 0 la_data_in[84]
port 272 nsew
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1750 90 0 0 la_data_in[85]
port 273 nsew
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1750 90 0 0 la_data_in[86]
port 274 nsew
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1750 90 0 0 la_data_in[87]
port 275 nsew
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1750 90 0 0 la_data_in[88]
port 276 nsew
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1750 90 0 0 la_data_in[89]
port 277 nsew
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1750 90 0 0 la_data_in[8]
port 278 nsew
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1750 90 0 0 la_data_in[90]
port 279 nsew
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1750 90 0 0 la_data_in[91]
port 280 nsew
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1750 90 0 0 la_data_in[92]
port 281 nsew
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1750 90 0 0 la_data_in[93]
port 282 nsew
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1750 90 0 0 la_data_in[94]
port 283 nsew
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1750 90 0 0 la_data_in[95]
port 284 nsew
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1750 90 0 0 la_data_in[96]
port 285 nsew
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1750 90 0 0 la_data_in[97]
port 286 nsew
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1750 90 0 0 la_data_in[98]
port 287 nsew
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1750 90 0 0 la_data_in[99]
port 288 nsew
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1750 90 0 0 la_data_in[9]
port 289 nsew
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1750 90 0 0 la_data_out[0]
port 290 nsew
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1750 90 0 0 la_data_out[100]
port 291 nsew
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1750 90 0 0 la_data_out[101]
port 292 nsew
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1750 90 0 0 la_data_out[102]
port 293 nsew
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1750 90 0 0 la_data_out[103]
port 294 nsew
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1750 90 0 0 la_data_out[104]
port 295 nsew
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1750 90 0 0 la_data_out[105]
port 296 nsew
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1750 90 0 0 la_data_out[106]
port 297 nsew
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1750 90 0 0 la_data_out[107]
port 298 nsew
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1750 90 0 0 la_data_out[108]
port 299 nsew
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1750 90 0 0 la_data_out[109]
port 300 nsew
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1750 90 0 0 la_data_out[10]
port 301 nsew
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1750 90 0 0 la_data_out[110]
port 302 nsew
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1750 90 0 0 la_data_out[111]
port 303 nsew
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1750 90 0 0 la_data_out[112]
port 304 nsew
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1750 90 0 0 la_data_out[113]
port 305 nsew
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1750 90 0 0 la_data_out[114]
port 306 nsew
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1750 90 0 0 la_data_out[115]
port 307 nsew
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1750 90 0 0 la_data_out[116]
port 308 nsew
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1750 90 0 0 la_data_out[117]
port 309 nsew
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1750 90 0 0 la_data_out[118]
port 310 nsew
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1750 90 0 0 la_data_out[119]
port 311 nsew
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1750 90 0 0 la_data_out[11]
port 312 nsew
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1750 90 0 0 la_data_out[120]
port 313 nsew
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1750 90 0 0 la_data_out[121]
port 314 nsew
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1750 90 0 0 la_data_out[122]
port 315 nsew
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1750 90 0 0 la_data_out[123]
port 316 nsew
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1750 90 0 0 la_data_out[124]
port 317 nsew
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1750 90 0 0 la_data_out[125]
port 318 nsew
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1750 90 0 0 la_data_out[126]
port 319 nsew
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1750 90 0 0 la_data_out[127]
port 320 nsew
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1750 90 0 0 la_data_out[12]
port 321 nsew
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1750 90 0 0 la_data_out[13]
port 322 nsew
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1750 90 0 0 la_data_out[14]
port 323 nsew
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1750 90 0 0 la_data_out[15]
port 324 nsew
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1750 90 0 0 la_data_out[16]
port 325 nsew
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1750 90 0 0 la_data_out[17]
port 326 nsew
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1750 90 0 0 la_data_out[18]
port 327 nsew
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1750 90 0 0 la_data_out[19]
port 328 nsew
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1750 90 0 0 la_data_out[1]
port 329 nsew
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1750 90 0 0 la_data_out[20]
port 330 nsew
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1750 90 0 0 la_data_out[21]
port 331 nsew
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1750 90 0 0 la_data_out[22]
port 332 nsew
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1750 90 0 0 la_data_out[23]
port 333 nsew
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1750 90 0 0 la_data_out[24]
port 334 nsew
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1750 90 0 0 la_data_out[25]
port 335 nsew
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1750 90 0 0 la_data_out[26]
port 336 nsew
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1750 90 0 0 la_data_out[27]
port 337 nsew
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1750 90 0 0 la_data_out[28]
port 338 nsew
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1750 90 0 0 la_data_out[29]
port 339 nsew
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1750 90 0 0 la_data_out[2]
port 340 nsew
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1750 90 0 0 la_data_out[30]
port 341 nsew
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1750 90 0 0 la_data_out[31]
port 342 nsew
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1750 90 0 0 la_data_out[32]
port 343 nsew
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1750 90 0 0 la_data_out[33]
port 344 nsew
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1750 90 0 0 la_data_out[34]
port 345 nsew
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1750 90 0 0 la_data_out[35]
port 346 nsew
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1750 90 0 0 la_data_out[36]
port 347 nsew
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1750 90 0 0 la_data_out[37]
port 348 nsew
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1750 90 0 0 la_data_out[38]
port 349 nsew
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1750 90 0 0 la_data_out[39]
port 350 nsew
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1750 90 0 0 la_data_out[3]
port 351 nsew
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1750 90 0 0 la_data_out[40]
port 352 nsew
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1750 90 0 0 la_data_out[41]
port 353 nsew
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1750 90 0 0 la_data_out[42]
port 354 nsew
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1750 90 0 0 la_data_out[43]
port 355 nsew
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1750 90 0 0 la_data_out[44]
port 356 nsew
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1750 90 0 0 la_data_out[45]
port 357 nsew
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1750 90 0 0 la_data_out[46]
port 358 nsew
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1750 90 0 0 la_data_out[47]
port 359 nsew
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1750 90 0 0 la_data_out[48]
port 360 nsew
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1750 90 0 0 la_data_out[49]
port 361 nsew
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1750 90 0 0 la_data_out[4]
port 362 nsew
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1750 90 0 0 la_data_out[50]
port 363 nsew
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1750 90 0 0 la_data_out[51]
port 364 nsew
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1750 90 0 0 la_data_out[52]
port 365 nsew
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1750 90 0 0 la_data_out[53]
port 366 nsew
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1750 90 0 0 la_data_out[54]
port 367 nsew
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1750 90 0 0 la_data_out[55]
port 368 nsew
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1750 90 0 0 la_data_out[56]
port 369 nsew
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1750 90 0 0 la_data_out[57]
port 370 nsew
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1750 90 0 0 la_data_out[58]
port 371 nsew
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1750 90 0 0 la_data_out[59]
port 372 nsew
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1750 90 0 0 la_data_out[5]
port 373 nsew
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1750 90 0 0 la_data_out[60]
port 374 nsew
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1750 90 0 0 la_data_out[61]
port 375 nsew
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1750 90 0 0 la_data_out[62]
port 376 nsew
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1750 90 0 0 la_data_out[63]
port 377 nsew
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1750 90 0 0 la_data_out[64]
port 378 nsew
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1750 90 0 0 la_data_out[65]
port 379 nsew
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1750 90 0 0 la_data_out[66]
port 380 nsew
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1750 90 0 0 la_data_out[67]
port 381 nsew
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1750 90 0 0 la_data_out[68]
port 382 nsew
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1750 90 0 0 la_data_out[69]
port 383 nsew
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1750 90 0 0 la_data_out[6]
port 384 nsew
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1750 90 0 0 la_data_out[70]
port 385 nsew
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1750 90 0 0 la_data_out[71]
port 386 nsew
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1750 90 0 0 la_data_out[72]
port 387 nsew
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1750 90 0 0 la_data_out[73]
port 388 nsew
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1750 90 0 0 la_data_out[74]
port 389 nsew
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1750 90 0 0 la_data_out[75]
port 390 nsew
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1750 90 0 0 la_data_out[76]
port 391 nsew
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1750 90 0 0 la_data_out[77]
port 392 nsew
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1750 90 0 0 la_data_out[78]
port 393 nsew
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1750 90 0 0 la_data_out[79]
port 394 nsew
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1750 90 0 0 la_data_out[7]
port 395 nsew
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1750 90 0 0 la_data_out[80]
port 396 nsew
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1750 90 0 0 la_data_out[81]
port 397 nsew
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1750 90 0 0 la_data_out[82]
port 398 nsew
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1750 90 0 0 la_data_out[83]
port 399 nsew
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1750 90 0 0 la_data_out[84]
port 400 nsew
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1750 90 0 0 la_data_out[85]
port 401 nsew
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1750 90 0 0 la_data_out[86]
port 402 nsew
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1750 90 0 0 la_data_out[87]
port 403 nsew
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1750 90 0 0 la_data_out[88]
port 404 nsew
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1750 90 0 0 la_data_out[89]
port 405 nsew
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1750 90 0 0 la_data_out[8]
port 406 nsew
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1750 90 0 0 la_data_out[90]
port 407 nsew
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1750 90 0 0 la_data_out[91]
port 408 nsew
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1750 90 0 0 la_data_out[92]
port 409 nsew
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1750 90 0 0 la_data_out[93]
port 410 nsew
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1750 90 0 0 la_data_out[94]
port 411 nsew
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1750 90 0 0 la_data_out[95]
port 412 nsew
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1750 90 0 0 la_data_out[96]
port 413 nsew
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1750 90 0 0 la_data_out[97]
port 414 nsew
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1750 90 0 0 la_data_out[98]
port 415 nsew
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1750 90 0 0 la_data_out[99]
port 416 nsew
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1750 90 0 0 la_data_out[9]
port 417 nsew
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1750 90 0 0 la_oenb[0]
port 418 nsew
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1750 90 0 0 la_oenb[100]
port 419 nsew
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1750 90 0 0 la_oenb[101]
port 420 nsew
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1750 90 0 0 la_oenb[102]
port 421 nsew
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1750 90 0 0 la_oenb[103]
port 422 nsew
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1750 90 0 0 la_oenb[104]
port 423 nsew
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1750 90 0 0 la_oenb[105]
port 424 nsew
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1750 90 0 0 la_oenb[106]
port 425 nsew
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1750 90 0 0 la_oenb[107]
port 426 nsew
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1750 90 0 0 la_oenb[108]
port 427 nsew
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1750 90 0 0 la_oenb[109]
port 428 nsew
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1750 90 0 0 la_oenb[10]
port 429 nsew
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1750 90 0 0 la_oenb[110]
port 430 nsew
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1750 90 0 0 la_oenb[111]
port 431 nsew
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1750 90 0 0 la_oenb[112]
port 432 nsew
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1750 90 0 0 la_oenb[113]
port 433 nsew
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1750 90 0 0 la_oenb[114]
port 434 nsew
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1750 90 0 0 la_oenb[115]
port 435 nsew
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1750 90 0 0 la_oenb[116]
port 436 nsew
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1750 90 0 0 la_oenb[117]
port 437 nsew
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1750 90 0 0 la_oenb[118]
port 438 nsew
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1750 90 0 0 la_oenb[119]
port 439 nsew
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1750 90 0 0 la_oenb[11]
port 440 nsew
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1750 90 0 0 la_oenb[120]
port 441 nsew
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1750 90 0 0 la_oenb[121]
port 442 nsew
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1750 90 0 0 la_oenb[122]
port 443 nsew
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1750 90 0 0 la_oenb[123]
port 444 nsew
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1750 90 0 0 la_oenb[124]
port 445 nsew
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1750 90 0 0 la_oenb[125]
port 446 nsew
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1750 90 0 0 la_oenb[126]
port 447 nsew
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1750 90 0 0 la_oenb[127]
port 448 nsew
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1750 90 0 0 la_oenb[12]
port 449 nsew
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1750 90 0 0 la_oenb[13]
port 450 nsew
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1750 90 0 0 la_oenb[14]
port 451 nsew
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1750 90 0 0 la_oenb[15]
port 452 nsew
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1750 90 0 0 la_oenb[16]
port 453 nsew
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1750 90 0 0 la_oenb[17]
port 454 nsew
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1750 90 0 0 la_oenb[18]
port 455 nsew
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1750 90 0 0 la_oenb[19]
port 456 nsew
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1750 90 0 0 la_oenb[1]
port 457 nsew
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1750 90 0 0 la_oenb[20]
port 458 nsew
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1750 90 0 0 la_oenb[21]
port 459 nsew
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1750 90 0 0 la_oenb[22]
port 460 nsew
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1750 90 0 0 la_oenb[23]
port 461 nsew
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1750 90 0 0 la_oenb[24]
port 462 nsew
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1750 90 0 0 la_oenb[25]
port 463 nsew
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1750 90 0 0 la_oenb[26]
port 464 nsew
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1750 90 0 0 la_oenb[27]
port 465 nsew
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1750 90 0 0 la_oenb[28]
port 466 nsew
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1750 90 0 0 la_oenb[29]
port 467 nsew
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1750 90 0 0 la_oenb[2]
port 468 nsew
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1750 90 0 0 la_oenb[30]
port 469 nsew
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1750 90 0 0 la_oenb[31]
port 470 nsew
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1750 90 0 0 la_oenb[32]
port 471 nsew
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1750 90 0 0 la_oenb[33]
port 472 nsew
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1750 90 0 0 la_oenb[34]
port 473 nsew
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1750 90 0 0 la_oenb[35]
port 474 nsew
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1750 90 0 0 la_oenb[36]
port 475 nsew
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1750 90 0 0 la_oenb[37]
port 476 nsew
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1750 90 0 0 la_oenb[38]
port 477 nsew
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1750 90 0 0 la_oenb[39]
port 478 nsew
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1750 90 0 0 la_oenb[3]
port 479 nsew
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1750 90 0 0 la_oenb[40]
port 480 nsew
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1750 90 0 0 la_oenb[41]
port 481 nsew
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1750 90 0 0 la_oenb[42]
port 482 nsew
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1750 90 0 0 la_oenb[43]
port 483 nsew
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1750 90 0 0 la_oenb[44]
port 484 nsew
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1750 90 0 0 la_oenb[45]
port 485 nsew
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1750 90 0 0 la_oenb[46]
port 486 nsew
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1750 90 0 0 la_oenb[47]
port 487 nsew
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1750 90 0 0 la_oenb[48]
port 488 nsew
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1750 90 0 0 la_oenb[49]
port 489 nsew
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1750 90 0 0 la_oenb[4]
port 490 nsew
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1750 90 0 0 la_oenb[50]
port 491 nsew
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1750 90 0 0 la_oenb[51]
port 492 nsew
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1750 90 0 0 la_oenb[52]
port 493 nsew
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1750 90 0 0 la_oenb[53]
port 494 nsew
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1750 90 0 0 la_oenb[54]
port 495 nsew
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1750 90 0 0 la_oenb[55]
port 496 nsew
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1750 90 0 0 la_oenb[56]
port 497 nsew
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1750 90 0 0 la_oenb[57]
port 498 nsew
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1750 90 0 0 la_oenb[58]
port 499 nsew
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1750 90 0 0 la_oenb[59]
port 500 nsew
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1750 90 0 0 la_oenb[5]
port 501 nsew
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1750 90 0 0 la_oenb[60]
port 502 nsew
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1750 90 0 0 la_oenb[61]
port 503 nsew
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1750 90 0 0 la_oenb[62]
port 504 nsew
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1750 90 0 0 la_oenb[63]
port 505 nsew
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1750 90 0 0 la_oenb[64]
port 506 nsew
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1750 90 0 0 la_oenb[65]
port 507 nsew
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1750 90 0 0 la_oenb[66]
port 508 nsew
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1750 90 0 0 la_oenb[67]
port 509 nsew
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1750 90 0 0 la_oenb[68]
port 510 nsew
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1750 90 0 0 la_oenb[69]
port 511 nsew
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1750 90 0 0 la_oenb[6]
port 512 nsew
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1750 90 0 0 la_oenb[70]
port 513 nsew
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1750 90 0 0 la_oenb[71]
port 514 nsew
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1750 90 0 0 la_oenb[72]
port 515 nsew
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1750 90 0 0 la_oenb[73]
port 516 nsew
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1750 90 0 0 la_oenb[74]
port 517 nsew
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1750 90 0 0 la_oenb[75]
port 518 nsew
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1750 90 0 0 la_oenb[76]
port 519 nsew
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1750 90 0 0 la_oenb[77]
port 520 nsew
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1750 90 0 0 la_oenb[78]
port 521 nsew
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1750 90 0 0 la_oenb[79]
port 522 nsew
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1750 90 0 0 la_oenb[7]
port 523 nsew
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1750 90 0 0 la_oenb[80]
port 524 nsew
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1750 90 0 0 la_oenb[81]
port 525 nsew
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1750 90 0 0 la_oenb[82]
port 526 nsew
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1750 90 0 0 la_oenb[83]
port 527 nsew
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1750 90 0 0 la_oenb[84]
port 528 nsew
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1750 90 0 0 la_oenb[85]
port 529 nsew
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1750 90 0 0 la_oenb[86]
port 530 nsew
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1750 90 0 0 la_oenb[87]
port 531 nsew
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1750 90 0 0 la_oenb[88]
port 532 nsew
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1750 90 0 0 la_oenb[89]
port 533 nsew
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1750 90 0 0 la_oenb[8]
port 534 nsew
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1750 90 0 0 la_oenb[90]
port 535 nsew
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1750 90 0 0 la_oenb[91]
port 536 nsew
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1750 90 0 0 la_oenb[92]
port 537 nsew
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1750 90 0 0 la_oenb[93]
port 538 nsew
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1750 90 0 0 la_oenb[94]
port 539 nsew
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1750 90 0 0 la_oenb[95]
port 540 nsew
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1750 90 0 0 la_oenb[96]
port 541 nsew
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1750 90 0 0 la_oenb[97]
port 542 nsew
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1750 90 0 0 la_oenb[98]
port 543 nsew
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1750 90 0 0 la_oenb[99]
port 544 nsew
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1750 90 0 0 la_oenb[9]
port 545 nsew
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1750 90 0 0 user_clock2
port 546 nsew
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1750 90 0 0 user_irq[0]
port 547 nsew
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1750 90 0 0 user_irq[1]
port 548 nsew
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1750 90 0 0 user_irq[2]
port 549 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1750 0 0 0 vccd1
port 550 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1750 0 0 0 vccd1
port 550 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1750 0 0 0 vccd2
port 551 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1750 0 0 0 vccd2
port 551 nsew
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1750 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1750 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1750 0 0 0 vdda1
port 552 nsew
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1750 0 0 0 vdda1
port 552 nsew
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1750 0 0 0 vdda2
port 553 nsew
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1750 0 0 0 vdda2
port 553 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 3000 180 0 0 vssa1
port 554 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 3000 180 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1750 0 0 0 vssa1
port 554 nsew
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1750 0 0 0 vssa1
port 554 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1750 0 0 0 vssa2
port 555 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1750 0 0 0 vssa2
port 555 nsew
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1750 0 0 0 vssd1
port 556 nsew
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1750 0 0 0 vssd1
port 556 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1750 0 0 0 vssd2
port 557 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1750 0 0 0 vssd2
port 557 nsew
flabel metal2 s 524 -800 636 480 0 FreeSans 1750 90 0 0 wb_clk_i
port 558 nsew
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1750 90 0 0 wb_rst_i
port 559 nsew
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1750 90 0 0 wbs_ack_o
port 560 nsew
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1750 90 0 0 wbs_adr_i[0]
port 561 nsew
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1750 90 0 0 wbs_adr_i[10]
port 562 nsew
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1750 90 0 0 wbs_adr_i[11]
port 563 nsew
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1750 90 0 0 wbs_adr_i[12]
port 564 nsew
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1750 90 0 0 wbs_adr_i[13]
port 565 nsew
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1750 90 0 0 wbs_adr_i[14]
port 566 nsew
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1750 90 0 0 wbs_adr_i[15]
port 567 nsew
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1750 90 0 0 wbs_adr_i[16]
port 568 nsew
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1750 90 0 0 wbs_adr_i[17]
port 569 nsew
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1750 90 0 0 wbs_adr_i[18]
port 570 nsew
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1750 90 0 0 wbs_adr_i[19]
port 571 nsew
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1750 90 0 0 wbs_adr_i[1]
port 572 nsew
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1750 90 0 0 wbs_adr_i[20]
port 573 nsew
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1750 90 0 0 wbs_adr_i[21]
port 574 nsew
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1750 90 0 0 wbs_adr_i[22]
port 575 nsew
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1750 90 0 0 wbs_adr_i[23]
port 576 nsew
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1750 90 0 0 wbs_adr_i[24]
port 577 nsew
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1750 90 0 0 wbs_adr_i[25]
port 578 nsew
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1750 90 0 0 wbs_adr_i[26]
port 579 nsew
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1750 90 0 0 wbs_adr_i[27]
port 580 nsew
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1750 90 0 0 wbs_adr_i[28]
port 581 nsew
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1750 90 0 0 wbs_adr_i[29]
port 582 nsew
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1750 90 0 0 wbs_adr_i[2]
port 583 nsew
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1750 90 0 0 wbs_adr_i[30]
port 584 nsew
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1750 90 0 0 wbs_adr_i[31]
port 585 nsew
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1750 90 0 0 wbs_adr_i[3]
port 586 nsew
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1750 90 0 0 wbs_adr_i[4]
port 587 nsew
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1750 90 0 0 wbs_adr_i[5]
port 588 nsew
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1750 90 0 0 wbs_adr_i[6]
port 589 nsew
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1750 90 0 0 wbs_adr_i[7]
port 590 nsew
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1750 90 0 0 wbs_adr_i[8]
port 591 nsew
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1750 90 0 0 wbs_adr_i[9]
port 592 nsew
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1750 90 0 0 wbs_cyc_i
port 593 nsew
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1750 90 0 0 wbs_dat_i[0]
port 594 nsew
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1750 90 0 0 wbs_dat_i[10]
port 595 nsew
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1750 90 0 0 wbs_dat_i[11]
port 596 nsew
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1750 90 0 0 wbs_dat_i[12]
port 597 nsew
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1750 90 0 0 wbs_dat_i[13]
port 598 nsew
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1750 90 0 0 wbs_dat_i[14]
port 599 nsew
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1750 90 0 0 wbs_dat_i[15]
port 600 nsew
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1750 90 0 0 wbs_dat_i[16]
port 601 nsew
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1750 90 0 0 wbs_dat_i[17]
port 602 nsew
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1750 90 0 0 wbs_dat_i[18]
port 603 nsew
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1750 90 0 0 wbs_dat_i[19]
port 604 nsew
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1750 90 0 0 wbs_dat_i[1]
port 605 nsew
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1750 90 0 0 wbs_dat_i[20]
port 606 nsew
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1750 90 0 0 wbs_dat_i[21]
port 607 nsew
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1750 90 0 0 wbs_dat_i[22]
port 608 nsew
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1750 90 0 0 wbs_dat_i[23]
port 609 nsew
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1750 90 0 0 wbs_dat_i[24]
port 610 nsew
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1750 90 0 0 wbs_dat_i[25]
port 611 nsew
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1750 90 0 0 wbs_dat_i[26]
port 612 nsew
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1750 90 0 0 wbs_dat_i[27]
port 613 nsew
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1750 90 0 0 wbs_dat_i[28]
port 614 nsew
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1750 90 0 0 wbs_dat_i[29]
port 615 nsew
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1750 90 0 0 wbs_dat_i[2]
port 616 nsew
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1750 90 0 0 wbs_dat_i[30]
port 617 nsew
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1750 90 0 0 wbs_dat_i[31]
port 618 nsew
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1750 90 0 0 wbs_dat_i[3]
port 619 nsew
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1750 90 0 0 wbs_dat_i[4]
port 620 nsew
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1750 90 0 0 wbs_dat_i[5]
port 621 nsew
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1750 90 0 0 wbs_dat_i[6]
port 622 nsew
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1750 90 0 0 wbs_dat_i[7]
port 623 nsew
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1750 90 0 0 wbs_dat_i[8]
port 624 nsew
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1750 90 0 0 wbs_dat_i[9]
port 625 nsew
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1750 90 0 0 wbs_dat_o[0]
port 626 nsew
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1750 90 0 0 wbs_dat_o[10]
port 627 nsew
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1750 90 0 0 wbs_dat_o[11]
port 628 nsew
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1750 90 0 0 wbs_dat_o[12]
port 629 nsew
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1750 90 0 0 wbs_dat_o[13]
port 630 nsew
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1750 90 0 0 wbs_dat_o[14]
port 631 nsew
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1750 90 0 0 wbs_dat_o[15]
port 632 nsew
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1750 90 0 0 wbs_dat_o[16]
port 633 nsew
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1750 90 0 0 wbs_dat_o[17]
port 634 nsew
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1750 90 0 0 wbs_dat_o[18]
port 635 nsew
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1750 90 0 0 wbs_dat_o[19]
port 636 nsew
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1750 90 0 0 wbs_dat_o[1]
port 637 nsew
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1750 90 0 0 wbs_dat_o[20]
port 638 nsew
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1750 90 0 0 wbs_dat_o[21]
port 639 nsew
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1750 90 0 0 wbs_dat_o[22]
port 640 nsew
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1750 90 0 0 wbs_dat_o[23]
port 641 nsew
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1750 90 0 0 wbs_dat_o[24]
port 642 nsew
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1750 90 0 0 wbs_dat_o[25]
port 643 nsew
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1750 90 0 0 wbs_dat_o[26]
port 644 nsew
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1750 90 0 0 wbs_dat_o[27]
port 645 nsew
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1750 90 0 0 wbs_dat_o[28]
port 646 nsew
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1750 90 0 0 wbs_dat_o[29]
port 647 nsew
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1750 90 0 0 wbs_dat_o[2]
port 648 nsew
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1750 90 0 0 wbs_dat_o[30]
port 649 nsew
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1750 90 0 0 wbs_dat_o[31]
port 650 nsew
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1750 90 0 0 wbs_dat_o[3]
port 651 nsew
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1750 90 0 0 wbs_dat_o[4]
port 652 nsew
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1750 90 0 0 wbs_dat_o[5]
port 653 nsew
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1750 90 0 0 wbs_dat_o[6]
port 654 nsew
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1750 90 0 0 wbs_dat_o[7]
port 655 nsew
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1750 90 0 0 wbs_dat_o[8]
port 656 nsew
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1750 90 0 0 wbs_dat_o[9]
port 657 nsew
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1750 90 0 0 wbs_sel_i[0]
port 658 nsew
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1750 90 0 0 wbs_sel_i[1]
port 659 nsew
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1750 90 0 0 wbs_sel_i[2]
port 660 nsew
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1750 90 0 0 wbs_sel_i[3]
port 661 nsew
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1750 90 0 0 wbs_stb_i
port 662 nsew
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1750 90 0 0 wbs_we_i
port 663 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

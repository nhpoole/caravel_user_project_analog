magic
tech sky130A
magscale 1 2
timestamp 1624134973
<< nwell >>
rect 10260 -57542 12494 -56702
<< pwell >>
rect 12118 -57600 12148 -57598
rect 12198 -57600 12410 -57598
rect 12118 -58256 12410 -57600
<< viali >>
rect 10342 -56772 10562 -56738
rect 11834 -56772 12036 -56738
rect 10294 -57408 10332 -56836
rect 12070 -57410 12106 -56834
rect 10342 -57506 10562 -57472
rect 11834 -57504 12036 -57470
rect 12238 -57586 12286 -57538
rect 12342 -57586 12390 -57538
rect 10366 -57708 10574 -57670
rect 11838 -57706 12036 -57668
rect 10294 -58124 10330 -57768
rect 12070 -58124 12108 -57768
rect 10364 -58220 10572 -58184
rect 11836 -58222 12038 -58186
<< metal1 >>
rect -74 -48 106 12
rect 53108 -40077 53114 -40017
rect 53174 -40077 53424 -40017
rect 30132 -41240 30192 -41148
rect 30132 -41306 30192 -41300
rect 30132 -41822 30192 -41816
rect 30132 -41888 30192 -41882
rect 57134 -41984 57194 -41978
rect 57034 -42044 57134 -41984
rect 57134 -42050 57194 -42044
rect 26980 -45164 26986 -45104
rect 27046 -45164 27052 -45104
rect 27774 -45164 27780 -45104
rect 27840 -45164 27846 -45104
rect 26980 -46920 26986 -46860
rect 27046 -46920 27052 -46860
rect 27774 -46920 27780 -46860
rect 27840 -46920 27846 -46860
rect 26980 -48434 26986 -48374
rect 27046 -48434 27052 -48374
rect 26976 -49676 26982 -49616
rect 27042 -49676 27048 -49616
rect 26980 -50912 26986 -50852
rect 27046 -50912 27052 -50852
rect 14762 -52948 14862 -52942
rect 27776 -53022 27782 -52962
rect 27842 -53022 27848 -52962
rect 14762 -53054 14862 -53048
rect 26374 -53624 26380 -53564
rect 26440 -53624 26446 -53564
rect 27774 -53624 27780 -53564
rect 27840 -53624 27846 -53564
rect 26380 -53734 26440 -53624
rect 14764 -53942 14864 -53936
rect 14764 -54048 14864 -54042
rect 14764 -54948 14864 -54942
rect 14764 -55054 14864 -55048
rect 27774 -55456 27780 -55396
rect 27840 -55456 27846 -55396
rect 10528 -56672 11876 -56612
rect 9350 -56724 9452 -56700
rect 9350 -57518 9372 -56724
rect 9436 -56726 10454 -56724
rect 10528 -56726 10588 -56672
rect 9436 -56738 10588 -56726
rect 9436 -56772 10342 -56738
rect 10562 -56772 10588 -56738
rect 9436 -56784 10588 -56772
rect 9436 -57094 9452 -56784
rect 10284 -56786 10588 -56784
rect 10284 -56836 10344 -56786
rect 10284 -57094 10294 -56836
rect 9436 -57154 10294 -57094
rect 9436 -57458 9452 -57154
rect 10284 -57408 10294 -57154
rect 10332 -57094 10344 -56836
rect 10394 -57094 10454 -56786
rect 10528 -56877 10588 -56786
rect 10784 -56720 10844 -56719
rect 11560 -56720 11620 -56714
rect 10784 -56780 11560 -56720
rect 10784 -56875 10844 -56780
rect 11042 -56877 11102 -56780
rect 11300 -56875 11360 -56780
rect 11560 -56875 11620 -56780
rect 11816 -56722 11876 -56672
rect 11816 -56738 12118 -56722
rect 11816 -56772 11834 -56738
rect 12036 -56772 12118 -56738
rect 11816 -56786 12118 -56772
rect 11816 -56877 11876 -56786
rect 10332 -57154 10454 -57094
rect 11944 -57092 12004 -56786
rect 12058 -56834 12118 -56786
rect 12058 -57092 12070 -56834
rect 11944 -57152 12070 -57092
rect 10332 -57408 10344 -57154
rect 10284 -57458 10344 -57408
rect 10396 -57458 10456 -57276
rect 10524 -57458 10584 -57370
rect 9436 -57472 10584 -57458
rect 9436 -57506 10342 -57472
rect 10562 -57506 10584 -57472
rect 9436 -57518 10584 -57506
rect 9350 -57536 9452 -57518
rect 10654 -57635 10714 -57265
rect 10912 -57486 10972 -57290
rect 10906 -57546 10912 -57486
rect 10972 -57546 10978 -57486
rect 10282 -57670 10586 -57660
rect 10282 -57708 10366 -57670
rect 10574 -57708 10586 -57670
rect 10648 -57695 10654 -57635
rect 10714 -57695 10720 -57635
rect 10282 -57720 10586 -57708
rect 10282 -57768 10342 -57720
rect 10282 -58124 10294 -57768
rect 10330 -58124 10342 -57768
rect 10396 -57908 10456 -57720
rect 10526 -57808 10586 -57720
rect 10654 -57895 10714 -57695
rect 10912 -57828 10972 -57546
rect 11170 -57635 11230 -57267
rect 11430 -57486 11490 -57272
rect 11424 -57546 11430 -57486
rect 11490 -57546 11496 -57486
rect 11164 -57695 11170 -57635
rect 11230 -57695 11236 -57635
rect 10912 -57894 10974 -57828
rect 10282 -58173 10342 -58124
rect 10398 -58173 10458 -57995
rect 10914 -58074 10974 -57894
rect 11170 -58014 11230 -57695
rect 11430 -58074 11490 -57546
rect 11688 -57635 11748 -57267
rect 11812 -57458 11872 -57370
rect 11946 -57458 12006 -57280
rect 12058 -57410 12070 -57152
rect 12106 -57210 12118 -56834
rect 15194 -56954 15562 -56894
rect 17356 -56954 17566 -56894
rect 12106 -57306 12184 -57210
rect 12106 -57410 12118 -57306
rect 12058 -57458 12118 -57410
rect 11812 -57470 12118 -57458
rect 11812 -57504 11834 -57470
rect 12036 -57504 12118 -57470
rect 11812 -57518 12118 -57504
rect 12176 -57532 12236 -57526
rect 12524 -57532 12584 -57526
rect 12236 -57538 12298 -57532
rect 12236 -57586 12238 -57538
rect 12286 -57586 12298 -57538
rect 12236 -57592 12298 -57586
rect 12330 -57538 12524 -57532
rect 12330 -57586 12342 -57538
rect 12390 -57586 12524 -57538
rect 12330 -57592 12524 -57586
rect 12176 -57598 12236 -57592
rect 12524 -57598 12584 -57592
rect 11688 -57897 11748 -57695
rect 11818 -57668 12120 -57658
rect 11818 -57706 11838 -57668
rect 12036 -57706 12120 -57668
rect 11818 -57718 12120 -57706
rect 11818 -57806 11878 -57718
rect 11946 -57904 12006 -57718
rect 12060 -57754 12120 -57718
rect 12060 -57768 12190 -57754
rect 10526 -58173 10586 -58084
rect 10282 -58184 10586 -58173
rect 10282 -58220 10364 -58184
rect 10572 -58220 10586 -58184
rect 10282 -58233 10586 -58220
rect 10282 -58390 10342 -58233
rect 10398 -58390 10458 -58233
rect 10526 -58390 10586 -58233
rect 10784 -58183 10844 -58083
rect 10908 -58134 10914 -58074
rect 10974 -58134 10980 -58074
rect 11044 -58183 11104 -58083
rect 11302 -58183 11362 -58085
rect 11424 -58134 11430 -58074
rect 11490 -58134 11496 -58074
rect 11558 -58183 11618 -58085
rect 11816 -58173 11876 -58082
rect 11944 -58173 12004 -58001
rect 12060 -58124 12070 -57768
rect 12108 -57850 12190 -57768
rect 12436 -57850 13132 -57754
rect 12108 -58124 12120 -57850
rect 12060 -58173 12120 -58124
rect 10784 -58243 11558 -58183
rect 11618 -58243 11624 -58183
rect 11816 -58186 12120 -58173
rect 11816 -58222 11836 -58186
rect 12038 -58222 12120 -58186
rect 11816 -58233 12120 -58222
rect 11816 -58390 11876 -58233
rect 11944 -58390 12004 -58233
rect 12060 -58390 12120 -58233
rect 10276 -58408 12130 -58390
rect 10276 -58514 10294 -58408
rect 12110 -58514 12130 -58408
rect 10276 -58528 12130 -58514
rect -3252 -72392 -3246 -72332
rect -3186 -72392 -3180 -72332
rect -2708 -72404 -2648 -71934
rect -2452 -72384 -2392 -71934
rect -28374 -72640 -28084 -72580
rect -24360 -72640 -24032 -72580
rect -20376 -72640 -20040 -72580
rect -16390 -72640 -16040 -72580
rect -12428 -72640 -12040 -72580
rect -8402 -72640 -8076 -72580
rect -392 -72640 -52 -72580
rect 3606 -72640 3958 -72580
rect -27092 -74870 -27032 -74054
rect -23092 -74868 -23032 -74034
rect -19092 -74868 -19032 -74042
rect -15092 -74868 -15032 -74048
rect -27098 -74930 -27092 -74870
rect -27032 -74930 -27026 -74870
rect -23098 -74928 -23092 -74868
rect -23032 -74928 -23026 -74868
rect -19098 -74928 -19092 -74868
rect -19032 -74928 -19026 -74868
rect -15098 -74928 -15092 -74868
rect -15032 -74928 -15026 -74868
rect -11092 -74870 -11032 -74034
rect -7092 -74870 -7032 -74036
rect -3092 -74868 -3032 -74034
rect 908 -74868 968 -74028
rect 4908 -74866 4968 -74040
rect -11098 -74930 -11092 -74870
rect -11032 -74930 -11026 -74870
rect -7098 -74930 -7092 -74870
rect -7032 -74930 -7026 -74870
rect -3098 -74928 -3092 -74868
rect -3032 -74928 -3026 -74868
rect 902 -74928 908 -74868
rect 968 -74928 974 -74868
rect 4902 -74926 4908 -74866
rect 4968 -74926 4974 -74866
<< via1 >>
rect 53114 -40077 53174 -40017
rect 30132 -41300 30192 -41240
rect 30132 -41882 30192 -41822
rect 57134 -42044 57194 -41984
rect 26986 -45164 27046 -45104
rect 27780 -45164 27840 -45104
rect 26986 -46920 27046 -46860
rect 27780 -46920 27840 -46860
rect 26986 -48434 27046 -48374
rect 26982 -49676 27042 -49616
rect 26986 -50912 27046 -50852
rect 14762 -53048 14862 -52948
rect 27782 -53022 27842 -52962
rect 26380 -53624 26440 -53564
rect 27780 -53624 27840 -53564
rect 14764 -54042 14864 -53942
rect 14764 -55048 14864 -54948
rect 27780 -55456 27840 -55396
rect 9372 -57518 9436 -56724
rect 11560 -56780 11620 -56720
rect 10912 -57546 10972 -57486
rect 10654 -57695 10714 -57635
rect 11430 -57546 11490 -57486
rect 11170 -57695 11230 -57635
rect 12176 -57592 12236 -57532
rect 12524 -57592 12584 -57532
rect 11688 -57695 11748 -57635
rect 10914 -58134 10974 -58074
rect 11430 -58134 11490 -58074
rect 11558 -58243 11618 -58183
rect 10294 -58514 12110 -58408
rect -3246 -72392 -3186 -72332
rect -27092 -74930 -27032 -74870
rect -23092 -74928 -23032 -74868
rect -19092 -74928 -19032 -74868
rect -15092 -74928 -15032 -74868
rect -11092 -74930 -11032 -74870
rect -7092 -74930 -7032 -74870
rect -3092 -74928 -3032 -74868
rect 908 -74928 968 -74868
rect 4908 -74926 4968 -74866
<< metal2 >>
rect 53114 -40017 53174 -40011
rect 52006 -40077 53114 -40017
rect 53114 -40083 53174 -40077
rect 49182 -41181 49191 -41091
rect 49281 -41181 49290 -41091
rect 51909 -41166 51918 -41106
rect 51978 -41166 53320 -41106
rect 30126 -41300 30132 -41240
rect 30192 -41300 30198 -41240
rect 30132 -41822 30192 -41300
rect 30126 -41882 30132 -41822
rect 30192 -41882 30198 -41822
rect 52380 -41962 52440 -41953
rect 52440 -42022 52500 -41962
rect 52380 -42031 52440 -42022
rect 57128 -42044 57134 -41984
rect 57194 -42044 57200 -41984
rect 58200 -41992 58452 -41932
rect 57134 -42132 57194 -42044
rect 57134 -42192 58450 -42132
rect 51994 -42542 53314 -42482
rect 53374 -42542 53383 -42482
rect 26986 -42942 27046 -42933
rect 26986 -43098 27046 -43002
rect 26986 -45104 27046 -45098
rect 27780 -45104 27840 -45098
rect 27046 -45164 27780 -45104
rect 26986 -45170 27046 -45164
rect 27780 -45170 27840 -45164
rect 26986 -46860 27046 -46854
rect 27780 -46860 27840 -46854
rect 27046 -46920 27780 -46860
rect 26986 -46926 27046 -46920
rect 27780 -46926 27840 -46920
rect 26986 -48374 27046 -48368
rect 27046 -48434 27900 -48374
rect 26986 -48440 27046 -48434
rect 26982 -49616 27042 -49610
rect 27042 -49676 28044 -49616
rect 26982 -49682 27042 -49676
rect 26986 -50852 27046 -50846
rect 27046 -50912 28070 -50852
rect 26986 -50918 27046 -50912
rect 14775 -51987 14865 -51978
rect 14775 -52086 14865 -52077
rect 14767 -52948 14857 -52944
rect 14756 -53048 14762 -52948
rect 14862 -53048 14868 -52948
rect 27782 -52962 27842 -52956
rect 26732 -53022 27782 -52962
rect 27782 -53028 27842 -53022
rect 14767 -53052 14857 -53048
rect 26380 -53564 26440 -53558
rect 27780 -53564 27840 -53558
rect 26440 -53624 27780 -53564
rect 26380 -53630 26440 -53624
rect 27780 -53630 27840 -53624
rect 14769 -53942 14859 -53938
rect 14758 -54042 14764 -53942
rect 14864 -54042 14870 -53942
rect 14769 -54046 14859 -54042
rect 14769 -54948 14859 -54944
rect 14758 -55048 14764 -54948
rect 14864 -55048 14870 -54948
rect 14769 -55052 14859 -55048
rect 27780 -55396 27840 -55390
rect 26320 -55456 27780 -55396
rect 27780 -55462 27840 -55456
rect 14779 -56339 14869 -56330
rect 14779 -56438 14869 -56429
rect 9350 -56724 9452 -56700
rect 9350 -57518 9372 -56724
rect 9436 -57518 9452 -56724
rect 11554 -56780 11560 -56720
rect 11620 -56780 12236 -56720
rect 9350 -57536 9452 -57518
rect 10912 -57486 10972 -57480
rect 11430 -57486 11490 -57480
rect 10972 -57546 11430 -57486
rect 12176 -57532 12236 -56780
rect 12524 -57532 12584 -57523
rect 10912 -57552 10972 -57546
rect 11430 -57552 11490 -57546
rect 12170 -57592 12176 -57532
rect 12236 -57592 12242 -57532
rect 12518 -57592 12524 -57532
rect 12584 -57592 12590 -57532
rect 12524 -57601 12584 -57592
rect 10654 -57635 10714 -57629
rect 11170 -57635 11230 -57629
rect 10643 -57695 10652 -57635
rect 10714 -57695 11170 -57635
rect 11230 -57695 11688 -57635
rect 11748 -57695 11754 -57635
rect 10654 -57701 10714 -57695
rect 11170 -57701 11230 -57695
rect 10914 -58074 10974 -58068
rect 10914 -58286 10974 -58134
rect 11430 -58074 11490 -58068
rect 11430 -58286 11490 -58134
rect 11558 -58183 11618 -58177
rect 11618 -58243 12526 -58183
rect 12586 -58243 12595 -58183
rect 11558 -58249 11618 -58243
rect 10914 -58346 13076 -58286
rect 10276 -58408 12130 -58390
rect 10276 -58514 10294 -58408
rect 12110 -58514 12130 -58408
rect 10276 -58528 12130 -58514
rect 13016 -59714 13076 -58346
rect 13007 -59774 13016 -59714
rect 13076 -59774 13085 -59714
rect -25067 -65195 -24977 -65186
rect -26400 -65274 -25067 -65214
rect -21031 -65197 -20941 -65188
rect -22446 -65274 -21031 -65214
rect -25067 -65294 -24977 -65285
rect -17109 -65197 -17019 -65188
rect -18454 -65274 -17109 -65214
rect -21031 -65296 -20941 -65287
rect -17109 -65296 -17019 -65287
rect -16087 -65197 -15997 -65188
rect -12623 -65197 -12533 -65188
rect -15997 -65274 -14694 -65214
rect -16087 -65296 -15997 -65287
rect -8033 -65199 -7943 -65190
rect -12533 -65274 -10656 -65214
rect -12623 -65296 -12533 -65287
rect -4097 -65197 -4007 -65188
rect -7943 -65274 -6710 -65214
rect -8033 -65298 -7943 -65289
rect -39 -65201 51 -65192
rect -4007 -65274 -2662 -65214
rect -4097 -65296 -4007 -65287
rect 4015 -65199 4105 -65190
rect 51 -65274 1320 -65214
rect -39 -65300 51 -65291
rect 4105 -65274 5342 -65214
rect 4015 -65298 4105 -65289
rect -26630 -65506 -26448 -65446
rect -26388 -65506 -26379 -65446
rect -22516 -65506 -22448 -65446
rect -22388 -65506 -22379 -65446
rect -18518 -65506 -18450 -65446
rect -18390 -65506 -18381 -65446
rect -14522 -65506 -14450 -65446
rect -14390 -65506 -14381 -65446
rect -10518 -65506 -10450 -65446
rect -10390 -65506 -10381 -65446
rect -6522 -65506 -6448 -65446
rect -6388 -65506 -6379 -65446
rect -2518 -65506 -2452 -65446
rect -2392 -65506 -2383 -65446
rect 1476 -65506 1552 -65446
rect 1612 -65506 1621 -65446
rect 5490 -65506 5554 -65446
rect 5614 -65506 5623 -65446
rect -26578 -67920 -26518 -67858
rect -22578 -67920 -22518 -67856
rect -18578 -67920 -18518 -67858
rect -14578 -67920 -14518 -67854
rect -10578 -67920 -10518 -67854
rect -6578 -67920 -6518 -67854
rect -2578 -67920 -2518 -67858
rect 1422 -67920 1482 -67854
rect -26587 -67980 -26578 -67920
rect -26518 -67980 -26509 -67920
rect -22587 -67980 -22578 -67920
rect -22518 -67980 -22509 -67920
rect -18587 -67980 -18578 -67920
rect -18518 -67980 -18509 -67920
rect -14587 -67980 -14578 -67920
rect -14518 -67980 -14509 -67920
rect -10587 -67980 -10578 -67920
rect -10518 -67980 -10509 -67920
rect -6587 -67980 -6578 -67920
rect -6518 -67980 -6509 -67920
rect -2587 -67980 -2578 -67920
rect -2518 -67980 -2509 -67920
rect 1413 -67980 1422 -67920
rect 1482 -67980 1491 -67920
rect 5422 -67922 5482 -67860
rect 5413 -67982 5422 -67922
rect 5482 -67982 5491 -67922
rect -26324 -69012 -25232 -68952
rect -25172 -69012 -25163 -68952
rect -22300 -69012 -21232 -68952
rect -21172 -69012 -21163 -68952
rect -18274 -69012 -17232 -68952
rect -17172 -69012 -17163 -68952
rect -14234 -69012 -13232 -68952
rect -13172 -69012 -13163 -68952
rect -10196 -69012 -9232 -68952
rect -9172 -69012 -9163 -68952
rect -6386 -69012 -5232 -68952
rect -5172 -69012 -5163 -68952
rect -2252 -69012 -1232 -68952
rect -1172 -69012 -1163 -68952
rect 1768 -69012 2768 -68952
rect 2828 -69012 2837 -68952
rect 5834 -69012 6768 -68952
rect 6828 -69012 6837 -68952
rect -25238 -72106 -25178 -72097
rect -21238 -72106 -21178 -72097
rect -17238 -72106 -17178 -72097
rect -13238 -72106 -13178 -72097
rect -9238 -72106 -9178 -72097
rect -5238 -72106 -5178 -72097
rect -1238 -72106 -1178 -72097
rect 2762 -72106 2822 -72097
rect 6762 -72106 6822 -72097
rect -26424 -72166 -25238 -72106
rect -22452 -72166 -21238 -72106
rect -18416 -72166 -17238 -72106
rect -14438 -72166 -13238 -72106
rect -10442 -72166 -9238 -72106
rect -6444 -72166 -5238 -72106
rect -2442 -72166 -1238 -72106
rect 1550 -72166 2762 -72106
rect 5566 -72166 6762 -72106
rect -25238 -72175 -25178 -72166
rect -21238 -72175 -21178 -72166
rect -17238 -72175 -17178 -72166
rect -13238 -72175 -13178 -72166
rect -9238 -72175 -9178 -72166
rect -5238 -72175 -5178 -72166
rect -1238 -72175 -1178 -72166
rect 2762 -72175 2822 -72166
rect 6762 -72175 6822 -72166
rect -3246 -72332 -3186 -72326
rect -3246 -72552 -3186 -72392
rect -27094 -72882 -27034 -72800
rect -23094 -72882 -23034 -72808
rect -19094 -72882 -19034 -72780
rect -15094 -72882 -15034 -72776
rect -11094 -72880 -11034 -72786
rect -27103 -72942 -27094 -72882
rect -27034 -72942 -27025 -72882
rect -23103 -72942 -23094 -72882
rect -23034 -72942 -23025 -72882
rect -19103 -72942 -19094 -72882
rect -19034 -72942 -19025 -72882
rect -15103 -72942 -15094 -72882
rect -15034 -72942 -15025 -72882
rect -11103 -72940 -11094 -72880
rect -11034 -72940 -11025 -72880
rect -7094 -72882 -7034 -72796
rect -3094 -72882 -3034 -72788
rect 906 -72882 966 -72786
rect -7103 -72942 -7094 -72882
rect -7034 -72942 -7025 -72882
rect -3103 -72942 -3094 -72882
rect -3034 -72942 -3025 -72882
rect 897 -72942 906 -72882
rect 966 -72942 975 -72882
rect 4897 -72942 4906 -72882
rect 4966 -72942 4975 -72882
rect -27092 -74870 -27032 -74864
rect -23092 -74868 -23032 -74862
rect -19092 -74868 -19032 -74862
rect -15092 -74868 -15032 -74862
rect -27101 -74930 -27092 -74870
rect -27032 -74930 -27023 -74870
rect -23101 -74928 -23092 -74868
rect -23032 -74928 -23023 -74868
rect -19101 -74928 -19092 -74868
rect -19032 -74928 -19023 -74868
rect -15101 -74928 -15092 -74868
rect -15032 -74928 -15023 -74868
rect -11092 -74870 -11032 -74864
rect -7092 -74870 -7032 -74864
rect -3092 -74868 -3032 -74862
rect 908 -74868 968 -74862
rect 4908 -74866 4968 -74860
rect -27092 -74936 -27032 -74930
rect -23092 -74934 -23032 -74928
rect -19092 -74934 -19032 -74928
rect -15092 -74934 -15032 -74928
rect -11101 -74930 -11092 -74870
rect -11032 -74930 -11023 -74870
rect -7101 -74930 -7092 -74870
rect -7032 -74930 -7023 -74870
rect -3101 -74928 -3092 -74868
rect -3032 -74928 -3023 -74868
rect 899 -74928 908 -74868
rect 968 -74928 977 -74868
rect 4899 -74926 4908 -74866
rect 4968 -74926 4977 -74866
rect -11092 -74936 -11032 -74930
rect -7092 -74936 -7032 -74930
rect -3092 -74934 -3032 -74928
rect 908 -74934 968 -74928
rect 4908 -74932 4968 -74926
<< via2 >>
rect 49191 -41181 49281 -41091
rect 51918 -41166 51978 -41106
rect 52380 -42022 52440 -41962
rect 53314 -42542 53374 -42482
rect 26986 -43002 27046 -42942
rect 14775 -52077 14865 -51987
rect 14767 -53043 14857 -52953
rect 14769 -54037 14859 -53947
rect 14769 -55043 14859 -54953
rect 14779 -56429 14869 -56339
rect 9372 -57518 9436 -56724
rect 12524 -57592 12584 -57532
rect 10652 -57695 10654 -57635
rect 10654 -57695 10712 -57635
rect 12526 -58243 12586 -58183
rect 10294 -58514 12110 -58408
rect 13016 -59774 13076 -59714
rect -25067 -65285 -24977 -65195
rect -21031 -65287 -20941 -65197
rect -17109 -65287 -17019 -65197
rect -16087 -65287 -15997 -65197
rect -12623 -65287 -12533 -65197
rect -8033 -65289 -7943 -65199
rect -4097 -65287 -4007 -65197
rect -39 -65291 51 -65201
rect 4015 -65289 4105 -65199
rect -26448 -65506 -26388 -65446
rect -22448 -65506 -22388 -65446
rect -18450 -65506 -18390 -65446
rect -14450 -65506 -14390 -65446
rect -10450 -65506 -10390 -65446
rect -6448 -65506 -6388 -65446
rect -2452 -65506 -2392 -65446
rect 1552 -65506 1612 -65446
rect 5554 -65506 5614 -65446
rect -26578 -67980 -26518 -67920
rect -22578 -67980 -22518 -67920
rect -18578 -67980 -18518 -67920
rect -14578 -67980 -14518 -67920
rect -10578 -67980 -10518 -67920
rect -6578 -67980 -6518 -67920
rect -2578 -67980 -2518 -67920
rect 1422 -67980 1482 -67920
rect 5422 -67982 5482 -67922
rect -25232 -69012 -25172 -68952
rect -21232 -69012 -21172 -68952
rect -17232 -69012 -17172 -68952
rect -13232 -69012 -13172 -68952
rect -9232 -69012 -9172 -68952
rect -5232 -69012 -5172 -68952
rect -1232 -69012 -1172 -68952
rect 2768 -69012 2828 -68952
rect 6768 -69012 6828 -68952
rect -25238 -72166 -25178 -72106
rect -21238 -72166 -21178 -72106
rect -17238 -72166 -17178 -72106
rect -13238 -72166 -13178 -72106
rect -9238 -72166 -9178 -72106
rect -5238 -72166 -5178 -72106
rect -1238 -72166 -1178 -72106
rect 2762 -72166 2822 -72106
rect 6762 -72166 6822 -72106
rect -27094 -72942 -27034 -72882
rect -23094 -72942 -23034 -72882
rect -19094 -72942 -19034 -72882
rect -15094 -72942 -15034 -72882
rect -11094 -72940 -11034 -72880
rect -7094 -72942 -7034 -72882
rect -3094 -72942 -3034 -72882
rect 906 -72942 966 -72882
rect 4906 -72942 4966 -72882
rect -27092 -74930 -27032 -74870
rect -23092 -74928 -23032 -74868
rect -19092 -74928 -19032 -74868
rect -15092 -74928 -15032 -74868
rect -11092 -74930 -11032 -74870
rect -7092 -74930 -7032 -74870
rect -3092 -74928 -3032 -74868
rect 908 -74928 968 -74868
rect 4908 -74926 4968 -74866
<< metal3 >>
rect -24278 -29944 -24178 -29206
rect -22172 -29944 -22072 -29206
rect -20066 -29944 -19966 -29206
rect -17960 -29944 -17860 -29206
rect -15854 -29944 -15754 -29206
rect -13748 -29944 -13648 -29206
rect -11642 -29944 -11542 -29206
rect -9536 -29944 -9436 -29206
rect -7430 -29944 -7330 -29206
rect -5324 -29944 -5224 -29206
rect -3218 -29944 -3118 -29206
rect -1112 -29944 -1012 -29206
rect 3060 -29944 3160 -29942
rect -26452 -30044 5328 -29944
rect -26392 -31934 -26292 -30782
rect -24286 -31934 -24178 -30044
rect -22172 -31934 -22072 -30044
rect -20066 -31934 -19966 -30044
rect -17960 -31934 -17860 -30044
rect -15854 -31934 -15754 -30044
rect -13748 -31934 -13648 -30044
rect -11642 -31934 -11542 -30044
rect -9536 -31934 -9436 -30044
rect -7430 -31934 -7330 -30044
rect -5324 -31934 -5224 -30044
rect -3218 -31934 -3118 -30044
rect -1112 -31934 -1012 -30044
rect 994 -31900 1094 -30044
rect 964 -31934 1094 -31900
rect 3060 -31934 3160 -30044
rect -26450 -31950 3160 -31934
rect 5228 -31950 5328 -30044
rect -26450 -32034 6076 -31950
rect -26392 -33956 -26292 -32034
rect -24286 -32806 -24178 -32034
rect -22172 -32408 -22072 -32034
rect -22172 -32806 -22034 -32408
rect -20066 -32806 -19936 -32034
rect -17960 -32806 -17792 -32034
rect -15854 -32806 -15754 -32034
rect -13748 -32806 -13648 -32034
rect -11642 -32806 -11542 -32034
rect -9536 -32806 -9436 -32034
rect -7430 -32806 -7330 -32034
rect -5324 -32806 -5224 -32034
rect -3218 -32806 -3118 -32034
rect -1112 -32362 -1012 -32034
rect -1134 -32806 -1012 -32362
rect 964 -32078 1094 -32034
rect 2355 -32050 6076 -32034
rect -24286 -33956 -24186 -32806
rect -22134 -33956 -22034 -32806
rect -20036 -33956 -19936 -32806
rect -17892 -33956 -17792 -32806
rect -26392 -34056 -17792 -33956
rect -26392 -35916 -26292 -34056
rect -24286 -35916 -24186 -34056
rect -22180 -35916 -22080 -34056
rect -26392 -36016 -22080 -35916
rect -20078 -35958 -19978 -35928
rect -15854 -35958 -15754 -33872
rect -13748 -33920 -13648 -33206
rect -11642 -33920 -11542 -33206
rect -9536 -33920 -9436 -33206
rect -7430 -33920 -7330 -33206
rect -5324 -33920 -5224 -33206
rect -15046 -34020 -3164 -33920
rect -13748 -35958 -13648 -34020
rect -11642 -35958 -11542 -34020
rect -9536 -35958 -9436 -34020
rect -7430 -35958 -7330 -34020
rect -5324 -35958 -5224 -34020
rect -3264 -35958 -3164 -34020
rect -1134 -33950 -1034 -32806
rect 964 -33950 1064 -32078
rect 3060 -33950 3160 -32050
rect 5228 -33950 5328 -32050
rect -1134 -34050 6076 -33950
rect 964 -35934 1064 -34050
rect 964 -35950 2978 -35934
rect 3060 -35950 3160 -34050
rect 5228 -35950 5328 -34050
rect -26392 -37942 -26292 -36016
rect -24286 -37942 -24186 -36016
rect -20134 -36058 -994 -35958
rect 964 -36034 6076 -35950
rect -26392 -38042 -24186 -37942
rect -22154 -37980 -22054 -37968
rect -20078 -37980 -19978 -36058
rect -13748 -36806 -13648 -36058
rect -11642 -36806 -11542 -36058
rect -9536 -36806 -9436 -36058
rect -7430 -36806 -7330 -36058
rect -5324 -36806 -5224 -36058
rect -26392 -39962 -26292 -38042
rect -24286 -39962 -24186 -38042
rect -22214 -38080 -19978 -37980
rect -26392 -40062 -24186 -39962
rect -22154 -39980 -22054 -38080
rect -20078 -39980 -19978 -38080
rect -17986 -38036 -3080 -37936
rect -17986 -39928 -17886 -38036
rect -15882 -39928 -15782 -38036
rect -26392 -41954 -26292 -40062
rect -24286 -41954 -24186 -40062
rect -22917 -40080 -19196 -39980
rect -17986 -40028 -15782 -39928
rect -12934 -40006 -7304 -39906
rect -26392 -42054 -24186 -41954
rect -22154 -41980 -22054 -40080
rect -20078 -41980 -19978 -40080
rect -26392 -43954 -26292 -42054
rect -24286 -43954 -24186 -42054
rect -22917 -42080 -19196 -41980
rect -27129 -44054 -23408 -43954
rect -22154 -43980 -22054 -42080
rect -20078 -43980 -19978 -42080
rect -26392 -45954 -26292 -44054
rect -24286 -45954 -24186 -44054
rect -22917 -44080 -19196 -43980
rect -27129 -46054 -23408 -45954
rect -22154 -45980 -22054 -44080
rect -20078 -45980 -19978 -44080
rect -26392 -47954 -26292 -46054
rect -24286 -47954 -24186 -46054
rect -22917 -46080 -19196 -45980
rect -27129 -48054 -23408 -47954
rect -22154 -47980 -22054 -46080
rect -20078 -47980 -19978 -46080
rect -26392 -49954 -26292 -48054
rect -24286 -49954 -24186 -48054
rect -22917 -48080 -19196 -47980
rect -27129 -50054 -23408 -49954
rect -22154 -49980 -22054 -48080
rect -20078 -49980 -19978 -48080
rect -17986 -49922 -17886 -40028
rect -13736 -40952 -13636 -40574
rect -15860 -41052 -13636 -40952
rect -7404 -40952 -7304 -40006
rect -5340 -39968 -5240 -38036
rect -3180 -39968 -3080 -38036
rect -5340 -40068 -3080 -39968
rect -15860 -48952 -15760 -41052
rect -13170 -41054 -7878 -40954
rect -7404 -41052 -5206 -40952
rect -13170 -41398 -13070 -41054
rect -7978 -41466 -7878 -41054
rect -10842 -42024 -9436 -41924
rect -14752 -42564 -14060 -42464
rect -14752 -47428 -14652 -42564
rect -11648 -42936 -11548 -42180
rect -13746 -43036 -11548 -42936
rect -9536 -42936 -9436 -42024
rect -6634 -42632 -6232 -42532
rect -9536 -43036 -7344 -42936
rect -13746 -46936 -13646 -43036
rect -10922 -44932 -10822 -44592
rect -10922 -45032 -10064 -44932
rect -10164 -45352 -10064 -45032
rect -7444 -46928 -7344 -43036
rect -13746 -47036 -11548 -46936
rect -14752 -47528 -14274 -47428
rect -11648 -47914 -11548 -47036
rect -9542 -47028 -7344 -46928
rect -9542 -47914 -9442 -47028
rect -6332 -47524 -6232 -42632
rect -6982 -47624 -6232 -47524
rect -11648 -48014 -9442 -47914
rect -13004 -48950 -12904 -48584
rect -9542 -48662 -9442 -48014
rect -8052 -48950 -7952 -48568
rect -5306 -48946 -5206 -41052
rect -15860 -49052 -13654 -48952
rect -13004 -49050 -7952 -48950
rect -7436 -49046 -5206 -48946
rect -13754 -49664 -13654 -49052
rect -7436 -49906 -7336 -49046
rect -26392 -51954 -26292 -50054
rect -24286 -51954 -24186 -50054
rect -22917 -50080 -19196 -49980
rect -17986 -50022 -15768 -49922
rect -14493 -50006 -6560 -49906
rect -3180 -49940 -3080 -40068
rect -1110 -39950 -1010 -36058
rect 964 -37918 1064 -36034
rect 2355 -36050 6076 -36034
rect 3060 -37918 3160 -36050
rect 964 -37950 3162 -37918
rect 5228 -37950 5328 -36050
rect 964 -38018 6076 -37950
rect 2355 -38050 6076 -38018
rect 3060 -39950 3160 -38050
rect 5228 -39950 5328 -38050
rect -1110 -40050 1110 -39950
rect 2355 -40050 6076 -39950
rect -1110 -41946 -1010 -40050
rect 1010 -41946 1110 -40050
rect -1154 -42046 1110 -41946
rect 3060 -41950 3160 -40050
rect 5228 -41950 5328 -40050
rect 49186 -41091 52004 -41086
rect 49186 -41181 49191 -41091
rect 49281 -41106 52004 -41091
rect 49281 -41166 51918 -41106
rect 51978 -41166 52004 -41106
rect 49281 -41181 52004 -41166
rect 49186 -41186 52004 -41181
rect -1110 -43916 -1010 -42046
rect 1010 -43916 1110 -42046
rect 2355 -42050 6076 -41950
rect 52310 -41962 52510 -41908
rect 52310 -42022 52380 -41962
rect 52440 -42022 52510 -41962
rect -1110 -44016 1110 -43916
rect 3060 -43950 3160 -42050
rect 5228 -43950 5328 -42050
rect 26958 -42937 27090 -42924
rect 26958 -43001 26981 -42937
rect 27051 -43001 27090 -42937
rect 26958 -43002 26986 -43001
rect 27046 -43002 27090 -43001
rect 26958 -43018 27090 -43002
rect -1110 -45948 -1010 -44016
rect 1010 -45948 1110 -44016
rect 2355 -44050 6076 -43950
rect -1154 -46048 1110 -45948
rect 3060 -45950 3160 -44050
rect 5228 -45950 5328 -44050
rect -1110 -47944 -1010 -46048
rect 1010 -47944 1110 -46048
rect 2355 -46050 6076 -45950
rect -1130 -48044 1110 -47944
rect 3060 -47950 3160 -46050
rect 5228 -47950 5328 -46050
rect -27129 -51956 -23408 -51954
rect -27129 -52054 -22126 -51956
rect -26392 -53954 -26292 -52054
rect -24286 -52056 -22126 -52054
rect -24286 -53954 -24186 -52056
rect -22226 -53954 -22126 -52056
rect -27129 -54054 -22080 -53954
rect -26392 -55954 -26292 -54054
rect -24286 -55954 -24186 -54054
rect -22180 -55954 -22080 -54054
rect -20078 -53970 -19978 -50080
rect -17986 -51980 -17886 -50022
rect -15868 -51980 -15768 -50022
rect -5324 -50040 -3080 -49940
rect -5324 -51980 -5224 -50040
rect -17986 -52080 -3918 -51980
rect -3180 -52114 -3080 -50040
rect -1110 -49926 -1010 -48044
rect 1010 -49926 1110 -48044
rect 2355 -48050 6076 -47950
rect -1110 -50026 1110 -49926
rect 3060 -49950 3160 -48050
rect 5228 -49950 5328 -48050
rect -1110 -51970 -1010 -50026
rect 1010 -51970 1110 -50026
rect 2355 -50050 6076 -49950
rect 3060 -51950 3160 -50050
rect 5228 -51950 5328 -50050
rect -1110 -52070 1110 -51970
rect 2355 -52050 6076 -51950
rect 7906 -51987 14870 -51982
rect -17970 -53970 -17870 -53966
rect -15864 -53970 -15764 -53206
rect -13758 -53970 -13658 -53206
rect -11652 -53970 -11552 -53206
rect -9546 -53970 -9446 -53206
rect -7440 -53970 -7340 -53206
rect -1110 -53970 -1010 -52070
rect 3060 -53950 3160 -52050
rect 5228 -53950 5328 -52050
rect 7906 -52077 14775 -51987
rect 14865 -52077 14870 -51987
rect 7906 -52082 14870 -52077
rect 8165 -52948 8263 -52943
rect 8164 -52949 14862 -52948
rect 8164 -53047 8165 -52949
rect 8263 -52953 14862 -52949
rect 8263 -53043 14767 -52953
rect 14857 -53043 14862 -52953
rect 8263 -53047 14862 -53043
rect 8164 -53048 14862 -53047
rect 8165 -53053 8263 -53048
rect 8138 -53947 14864 -53942
rect -20078 -54070 -1010 -53970
rect 1010 -54050 6076 -53950
rect 8138 -54037 14769 -53947
rect 14859 -54037 14864 -53947
rect 8138 -54042 14864 -54037
rect -27129 -56054 -19912 -55954
rect -26392 -57954 -26292 -56054
rect -24286 -57930 -24186 -56054
rect -22156 -57930 -22056 -56054
rect -20012 -57206 -19912 -56054
rect -17970 -55976 -17870 -54070
rect -15864 -55976 -15764 -54070
rect -13758 -55976 -13658 -54070
rect -11652 -55976 -11552 -54070
rect -9546 -55976 -9446 -54070
rect -7440 -55976 -7340 -54070
rect -5340 -55976 -5240 -54070
rect 1010 -55950 1110 -54050
rect 3060 -55950 3160 -54050
rect 5228 -55950 5328 -54050
rect 8163 -54948 8261 -54943
rect 8162 -54949 14864 -54948
rect 8162 -55047 8163 -54949
rect 8261 -54953 14864 -54949
rect 8261 -55043 14769 -54953
rect 14859 -55043 14864 -54953
rect 8261 -55047 14864 -55043
rect 8162 -55048 14864 -55047
rect 8163 -55053 8261 -55048
rect -17970 -56076 -5240 -55976
rect -3278 -56050 5328 -55950
rect -15864 -56806 -15764 -56076
rect -13758 -56806 -13658 -56076
rect -11652 -56806 -11552 -56076
rect -9546 -56806 -9446 -56076
rect -7440 -56806 -7340 -56076
rect -3278 -57206 -3178 -56050
rect -1156 -57206 -1056 -56050
rect 1010 -57206 1110 -56050
rect -20060 -57930 -19912 -57206
rect -17954 -57930 -17854 -57206
rect -15848 -57930 -15748 -57206
rect -13742 -57930 -13642 -57206
rect -11636 -57930 -11536 -57206
rect -9530 -57930 -9430 -57206
rect -7424 -57930 -7324 -57206
rect -5318 -57930 -5218 -57206
rect -3278 -57930 -3112 -57206
rect -1156 -57930 -1006 -57206
rect 1000 -57930 1110 -57206
rect 3060 -57206 3160 -56050
rect 3060 -57930 3206 -57206
rect 5228 -57930 5328 -56050
rect 8100 -56339 14874 -56334
rect 8100 -56429 14779 -56339
rect 14869 -56429 14874 -56339
rect 8100 -56434 14874 -56429
rect 9350 -56724 9452 -56700
rect 9350 -57518 9372 -56724
rect 9436 -57518 9452 -56724
rect 9350 -57536 9452 -57518
rect 12504 -57532 12604 -57512
rect 12504 -57592 12524 -57532
rect 12584 -57592 12604 -57532
rect 8086 -57635 10734 -57614
rect 8086 -57695 10652 -57635
rect 10712 -57695 10734 -57635
rect 8086 -57712 10734 -57695
rect 8086 -57714 10652 -57712
rect -24286 -57954 5328 -57930
rect -27129 -58030 5328 -57954
rect -27129 -58054 -23408 -58030
rect -26392 -59206 -26292 -58054
rect -26392 -60076 -26344 -59206
rect -24286 -59946 -24186 -58054
rect -22166 -58072 -22056 -58030
rect -20060 -58072 -19912 -58030
rect -22166 -59946 -22066 -58072
rect -20060 -59946 -19960 -58072
rect -17954 -59946 -17854 -58030
rect -15848 -59946 -15748 -58030
rect -13742 -59946 -13642 -58030
rect -11636 -59946 -11536 -58030
rect -9530 -59946 -9430 -58030
rect -7424 -59946 -7324 -58030
rect -5318 -59946 -5218 -58030
rect -3278 -58050 -3112 -58030
rect -3212 -59946 -3112 -58050
rect -1156 -58118 -1006 -58030
rect -1106 -59946 -1006 -58118
rect 1000 -58142 1110 -58030
rect 1000 -59946 1100 -58142
rect 3106 -59946 3206 -58030
rect 5228 -59946 5328 -58030
rect 12504 -58183 12604 -57592
rect 12504 -58243 12526 -58183
rect 12586 -58243 12604 -58183
rect 10276 -58408 12130 -58390
rect 10276 -58514 10294 -58408
rect 12110 -58514 12130 -58408
rect 10276 -58528 12130 -58514
rect -26244 -60046 5328 -59946
rect -25270 -63286 -25170 -60046
rect -24286 -60066 -24186 -60046
rect -22166 -60114 -22066 -60046
rect -20060 -60806 -19960 -60046
rect -17954 -60806 -17854 -60046
rect -15848 -60806 -15748 -60046
rect -13742 -60806 -13642 -60046
rect -11636 -60806 -11536 -60046
rect -9530 -60806 -9430 -60046
rect -7424 -60806 -7324 -60046
rect -5318 -60806 -5218 -60046
rect -3212 -60806 -3112 -60046
rect -1106 -60806 -1006 -60046
rect 1000 -60806 1100 -60046
rect 3106 -60806 3206 -60046
rect -9938 -63001 -9838 -63000
rect -14752 -63009 -14652 -63008
rect -16848 -63011 -16748 -63010
rect -18964 -63015 -18864 -63014
rect -18969 -63113 -18963 -63015
rect -18865 -63113 -18859 -63015
rect -16853 -63109 -16847 -63011
rect -16749 -63109 -16743 -63011
rect -14757 -63107 -14751 -63009
rect -14653 -63107 -14647 -63009
rect -10592 -63011 -10492 -63010
rect -12628 -63019 -12528 -63018
rect -25270 -63386 -24972 -63286
rect -18964 -63326 -18864 -63113
rect -16848 -63310 -16748 -63109
rect -25072 -65195 -24972 -63386
rect -25072 -65285 -25067 -65195
rect -24977 -65285 -24972 -65195
rect -25072 -65290 -24972 -65285
rect -21036 -63426 -18864 -63326
rect -17114 -63410 -16748 -63310
rect -21036 -65197 -20936 -63426
rect -21036 -65287 -21031 -65197
rect -20941 -65287 -20936 -65197
rect -21036 -65292 -20936 -65287
rect -17114 -65197 -17014 -63410
rect -14752 -63634 -14652 -63107
rect -12633 -63117 -12627 -63019
rect -12529 -63117 -12523 -63019
rect -10597 -63109 -10591 -63011
rect -10493 -63109 -10487 -63011
rect -9943 -63099 -9937 -63001
rect -9839 -63099 -9833 -63001
rect -8496 -63019 -8396 -63018
rect -17114 -65287 -17109 -65197
rect -17019 -65287 -17014 -65197
rect -17114 -65292 -17014 -65287
rect -16092 -63734 -14652 -63634
rect -16092 -65197 -15992 -63734
rect -16092 -65287 -16087 -65197
rect -15997 -65287 -15992 -65197
rect -16092 -65292 -15992 -65287
rect -12628 -65197 -12528 -63117
rect -10592 -64004 -10492 -63109
rect -9938 -63640 -9838 -63099
rect -8501 -63117 -8495 -63019
rect -8397 -63117 -8391 -63019
rect -7927 -63022 -7829 -63017
rect -7928 -63023 4110 -63022
rect -8496 -63322 -8396 -63117
rect -7928 -63121 -7927 -63023
rect -7829 -63121 4110 -63023
rect -7928 -63122 4110 -63121
rect -7927 -63127 -7829 -63122
rect -8496 -63422 56 -63322
rect -9938 -63740 -4002 -63640
rect -10592 -64104 -7938 -64004
rect -12628 -65287 -12623 -65197
rect -12533 -65287 -12528 -65197
rect -12628 -65292 -12528 -65287
rect -8038 -65199 -7938 -64104
rect -8038 -65289 -8033 -65199
rect -7943 -65289 -7938 -65199
rect -8038 -65294 -7938 -65289
rect -4102 -65197 -4002 -63740
rect -4102 -65287 -4097 -65197
rect -4007 -65287 -4002 -65197
rect -4102 -65292 -4002 -65287
rect -44 -65201 56 -63422
rect -44 -65291 -39 -65201
rect 51 -65291 56 -65201
rect -44 -65296 56 -65291
rect 4010 -65199 4110 -63122
rect 4010 -65289 4015 -65199
rect 4105 -65289 4110 -65199
rect 4010 -65294 4110 -65289
rect 12504 -65426 12604 -58243
rect 52310 -59666 52510 -42022
rect 53309 -42482 53379 -42477
rect 53309 -42542 53314 -42482
rect 53374 -42542 53379 -42482
rect 53309 -42547 53379 -42542
rect -26472 -65446 12604 -65426
rect -26472 -65506 -26448 -65446
rect -26388 -65506 -22448 -65446
rect -22388 -65506 -18450 -65446
rect -18390 -65506 -14450 -65446
rect -14390 -65506 -10450 -65446
rect -10390 -65506 -6448 -65446
rect -6388 -65506 -2452 -65446
rect -2392 -65506 1552 -65446
rect 1612 -65506 5554 -65446
rect 5614 -65506 12604 -65446
rect -26472 -65526 12604 -65506
rect 12962 -59714 52510 -59666
rect 12962 -59774 13016 -59714
rect 13076 -59774 52510 -59714
rect 12962 -59866 52510 -59774
rect -28296 -67920 5506 -67902
rect -28296 -67980 -26578 -67920
rect -26518 -67980 -22578 -67920
rect -22518 -67980 -18578 -67920
rect -18518 -67980 -14578 -67920
rect -14518 -67980 -10578 -67920
rect -10518 -67980 -6578 -67920
rect -6518 -67980 -2578 -67920
rect -2518 -67980 1422 -67920
rect 1482 -67922 5506 -67920
rect 1482 -67980 5422 -67922
rect -28296 -67982 5422 -67980
rect 5482 -67982 5506 -67922
rect -28296 -68002 5506 -67982
rect -25254 -68952 -25154 -68924
rect -25254 -69012 -25232 -68952
rect -25172 -69012 -25154 -68952
rect -25254 -72106 -25154 -69012
rect -25254 -72166 -25238 -72106
rect -25178 -72166 -25154 -72106
rect -25254 -72192 -25154 -72166
rect -21254 -68952 -21154 -68924
rect -21254 -69012 -21232 -68952
rect -21172 -69012 -21154 -68952
rect -21254 -72106 -21154 -69012
rect -21254 -72166 -21238 -72106
rect -21178 -72166 -21154 -72106
rect -21254 -72192 -21154 -72166
rect -17254 -68952 -17154 -68924
rect -17254 -69012 -17232 -68952
rect -17172 -69012 -17154 -68952
rect -17254 -72106 -17154 -69012
rect -17254 -72166 -17238 -72106
rect -17178 -72166 -17154 -72106
rect -17254 -72192 -17154 -72166
rect -13254 -68952 -13154 -68924
rect -13254 -69012 -13232 -68952
rect -13172 -69012 -13154 -68952
rect -13254 -72106 -13154 -69012
rect -13254 -72166 -13238 -72106
rect -13178 -72166 -13154 -72106
rect -13254 -72192 -13154 -72166
rect -9254 -68952 -9154 -68924
rect -9254 -69012 -9232 -68952
rect -9172 -69012 -9154 -68952
rect -9254 -72106 -9154 -69012
rect -9254 -72166 -9238 -72106
rect -9178 -72166 -9154 -72106
rect -9254 -72192 -9154 -72166
rect -5254 -68952 -5154 -68924
rect -5254 -69012 -5232 -68952
rect -5172 -69012 -5154 -68952
rect -5254 -72106 -5154 -69012
rect -5254 -72166 -5238 -72106
rect -5178 -72166 -5154 -72106
rect -5254 -72192 -5154 -72166
rect -1254 -68952 -1154 -68924
rect -1254 -69012 -1232 -68952
rect -1172 -69012 -1154 -68952
rect -1254 -72106 -1154 -69012
rect -1254 -72166 -1238 -72106
rect -1178 -72166 -1154 -72106
rect -1254 -72192 -1154 -72166
rect 2746 -68952 2846 -68924
rect 2746 -69012 2768 -68952
rect 2828 -69012 2846 -68952
rect 2746 -72106 2846 -69012
rect 2746 -72166 2762 -72106
rect 2822 -72166 2846 -72106
rect 2746 -72192 2846 -72166
rect 6746 -68952 6846 -68924
rect 6746 -69012 6768 -68952
rect 6828 -69012 6846 -68952
rect 6746 -72106 6846 -69012
rect 6746 -72166 6762 -72106
rect 6822 -72166 6846 -72106
rect 6746 -72192 6846 -72166
rect 12962 -72808 13162 -59866
rect 4844 -72864 13162 -72808
rect -28500 -72880 13162 -72864
rect -28500 -72882 -11094 -72880
rect -28500 -72942 -27094 -72882
rect -27034 -72942 -23094 -72882
rect -23034 -72942 -19094 -72882
rect -19034 -72942 -15094 -72882
rect -15034 -72940 -11094 -72882
rect -11034 -72882 13162 -72880
rect -11034 -72940 -7094 -72882
rect -15034 -72942 -7094 -72940
rect -7034 -72942 -3094 -72882
rect -3034 -72942 906 -72882
rect 966 -72942 4906 -72882
rect 4966 -72942 13162 -72882
rect -28500 -72964 13162 -72942
rect 4844 -73008 13162 -72964
rect -28238 -74866 4986 -74848
rect -28238 -74868 4908 -74866
rect -28238 -74870 -23092 -74868
rect -28238 -74930 -27092 -74870
rect -27032 -74928 -23092 -74870
rect -23032 -74928 -19092 -74868
rect -19032 -74928 -15092 -74868
rect -15032 -74870 -3092 -74868
rect -15032 -74928 -11092 -74870
rect -27032 -74930 -11092 -74928
rect -11032 -74930 -7092 -74870
rect -7032 -74928 -3092 -74870
rect -3032 -74928 908 -74868
rect 968 -74926 4908 -74868
rect 4968 -74926 4986 -74866
rect 968 -74928 4986 -74926
rect -7032 -74930 4986 -74928
rect -28238 -74948 4986 -74930
<< via3 >>
rect 26981 -42942 27051 -42937
rect 26981 -43001 26986 -42942
rect 26986 -43001 27046 -42942
rect 27046 -43001 27051 -42942
rect 8165 -53047 8263 -52949
rect 8163 -55047 8261 -54949
rect 9372 -57518 9436 -56724
rect 10294 -58514 12110 -58408
rect -18963 -63113 -18865 -63015
rect -16847 -63109 -16749 -63011
rect -14751 -63107 -14653 -63009
rect -12627 -63117 -12529 -63019
rect -10591 -63109 -10493 -63011
rect -9937 -63099 -9839 -63001
rect -8495 -63117 -8397 -63019
rect -7927 -63121 -7829 -63023
<< metal4 >>
rect 7330 -27958 8260 -27942
rect -28478 -28058 8276 -27958
rect -28470 -28948 -28370 -28058
rect -27640 -28948 -27540 -28058
rect -26348 -28948 -26248 -28058
rect -24242 -28948 -24142 -28058
rect -22136 -28948 -22036 -28058
rect -20030 -28948 -19930 -28058
rect -17924 -28948 -17824 -28058
rect -15818 -28948 -15718 -28058
rect -13712 -28948 -13612 -28058
rect -11606 -28948 -11506 -28058
rect -9500 -28948 -9400 -28058
rect -7394 -28948 -7294 -28058
rect -5288 -28948 -5188 -28058
rect -3182 -28948 -3082 -28058
rect -1076 -28948 -976 -28058
rect 1030 -28948 1130 -28058
rect 3136 -28948 3236 -28058
rect 5242 -28948 5342 -28058
rect 7368 -28948 7468 -28058
rect 8160 -28948 8260 -28058
rect 9588 -28378 11212 -27578
rect 48760 -28378 50552 -27578
rect -28470 -29048 8260 -28948
rect -28470 -29938 -28370 -29048
rect -27640 -29938 -27540 -29048
rect -28470 -30038 -27540 -29938
rect -28470 -30948 -28370 -30038
rect -27640 -30948 -27540 -30038
rect -26348 -30948 -26248 -29048
rect -24242 -30948 -24142 -29048
rect -22136 -30948 -22036 -29048
rect -20030 -30948 -19930 -29048
rect -17924 -30948 -17824 -29048
rect -15818 -30948 -15718 -29048
rect -13712 -30948 -13612 -29048
rect -11606 -30948 -11506 -29048
rect -9500 -30948 -9400 -29048
rect -7394 -30948 -7294 -29048
rect -5288 -30948 -5188 -29048
rect -3182 -30948 -3082 -29048
rect -1076 -30948 -976 -29048
rect 1030 -30948 1130 -29048
rect 3136 -30948 3236 -29048
rect 5242 -30948 5342 -29048
rect 7368 -29942 7468 -29048
rect 8160 -29942 8260 -29048
rect 7330 -30042 8260 -29942
rect 7368 -30948 7468 -30042
rect 8160 -30948 8260 -30042
rect -28470 -31048 8260 -30948
rect -28470 -31938 -28370 -31048
rect -27640 -31938 -27540 -31048
rect -28470 -32038 -27540 -31938
rect -28470 -32948 -28370 -32038
rect -27640 -32948 -27540 -32038
rect -26348 -32948 -26248 -31048
rect -24242 -32948 -24142 -31048
rect -22136 -32948 -22036 -31048
rect -20030 -32948 -19930 -31048
rect -17924 -32948 -17824 -31048
rect -15818 -32948 -15718 -31048
rect -13712 -32948 -13612 -31048
rect -11606 -32948 -11506 -31048
rect -9500 -32948 -9400 -31048
rect -7394 -32948 -7294 -31048
rect -5288 -32948 -5188 -31048
rect -3182 -32948 -3082 -31048
rect -1076 -32948 -976 -31048
rect 1030 -32948 1130 -31048
rect 3136 -32948 3236 -31048
rect 5242 -32948 5342 -31048
rect 7368 -31942 7468 -31048
rect 8160 -31942 8260 -31048
rect 7330 -32042 8260 -31942
rect 7368 -32948 7468 -32042
rect 8160 -32948 8260 -32042
rect -28470 -33048 8260 -32948
rect -28470 -33938 -28370 -33048
rect -27640 -33938 -27540 -33048
rect -28470 -34038 -27540 -33938
rect -28470 -34948 -28370 -34038
rect -27640 -34948 -27540 -34038
rect -26348 -34948 -26248 -33048
rect -24242 -34948 -24142 -33048
rect -22136 -34948 -22036 -33048
rect -20030 -34948 -19930 -33048
rect -17924 -34948 -17824 -33048
rect -15818 -34948 -15718 -33048
rect -13712 -34948 -13612 -33048
rect -11606 -34948 -11506 -33048
rect -9500 -34948 -9400 -33048
rect -7394 -34948 -7294 -33048
rect -5288 -34948 -5188 -33048
rect -3182 -34948 -3082 -33048
rect -1076 -34948 -976 -33048
rect 1030 -34948 1130 -33048
rect 3136 -34948 3236 -33048
rect 5242 -34948 5342 -33048
rect 7368 -33942 7468 -33048
rect 8160 -33942 8260 -33048
rect 7330 -34042 8260 -33942
rect 7368 -34948 7468 -34042
rect 8160 -34948 8260 -34042
rect -28470 -35048 8260 -34948
rect -28470 -35938 -28370 -35048
rect -27640 -35938 -27540 -35048
rect -28470 -36038 -27540 -35938
rect -28470 -36948 -28370 -36038
rect -27640 -36948 -27540 -36038
rect -26348 -36948 -26248 -35048
rect -24242 -36948 -24142 -35048
rect -22136 -36948 -22036 -35048
rect -20030 -36948 -19930 -35048
rect -17924 -36948 -17824 -35048
rect -15818 -36948 -15718 -35048
rect -13712 -36948 -13612 -35048
rect -11606 -36948 -11506 -35048
rect -9500 -36948 -9400 -35048
rect -7394 -36948 -7294 -35048
rect -5288 -36948 -5188 -35048
rect -3182 -36948 -3082 -35048
rect -1076 -36948 -976 -35048
rect 1030 -36948 1130 -35048
rect 3136 -36948 3236 -35048
rect 5242 -36948 5342 -35048
rect 7368 -35942 7468 -35048
rect 8160 -35942 8260 -35048
rect 7330 -36042 8260 -35942
rect 7368 -36948 7468 -36042
rect 8160 -36948 8260 -36042
rect -28470 -37048 8260 -36948
rect -28470 -37938 -28370 -37048
rect -27640 -37938 -27540 -37048
rect -28470 -38038 -27540 -37938
rect -28470 -38948 -28370 -38038
rect -27640 -38948 -27540 -38038
rect -26348 -38948 -26248 -37048
rect -24242 -38948 -24142 -37048
rect -22136 -38948 -22036 -37048
rect -20030 -38948 -19930 -37048
rect -17924 -38948 -17824 -37048
rect -15818 -38948 -15718 -37048
rect -13712 -38948 -13612 -37048
rect -11606 -38948 -11506 -37048
rect -9500 -38948 -9400 -37048
rect -7394 -38948 -7294 -37048
rect -5288 -38948 -5188 -37048
rect -3182 -38948 -3082 -37048
rect -1076 -38948 -976 -37048
rect 1030 -38948 1130 -37048
rect 3136 -38948 3236 -37048
rect 5242 -38948 5342 -37048
rect 7368 -37942 7468 -37048
rect 8160 -37942 8260 -37048
rect 7330 -38042 8260 -37942
rect 7368 -38948 7468 -38042
rect 8160 -38948 8260 -38042
rect -28470 -39048 8260 -38948
rect -28470 -39938 -28370 -39048
rect -27640 -39938 -27540 -39048
rect -28470 -40038 -27540 -39938
rect -28470 -40948 -28370 -40038
rect -27640 -40948 -27540 -40038
rect -26348 -40948 -26248 -39048
rect -24242 -40948 -24142 -39048
rect -22136 -40948 -22036 -39048
rect -20030 -40948 -19930 -39048
rect -17924 -40948 -17824 -39048
rect -15818 -40948 -15718 -39048
rect -13712 -40948 -13612 -39048
rect -11606 -40948 -11506 -39048
rect -9500 -40948 -9400 -39048
rect -7394 -40948 -7294 -39048
rect -5288 -40948 -5188 -39048
rect -3182 -40948 -3082 -39048
rect -1076 -40948 -976 -39048
rect 1030 -40948 1130 -39048
rect 3136 -40948 3236 -39048
rect 5242 -40948 5342 -39048
rect 7368 -39942 7468 -39048
rect 8160 -39942 8260 -39048
rect 50552 -38704 52664 -38680
rect 50552 -39456 50576 -38704
rect 51328 -39456 52664 -38704
rect 50552 -39480 52664 -39456
rect 7330 -40042 8260 -39942
rect 7368 -40948 7468 -40042
rect 8160 -40948 8260 -40042
rect -28470 -41048 8260 -40948
rect -28470 -41938 -28370 -41048
rect -27640 -41938 -27540 -41048
rect -28470 -42038 -27540 -41938
rect -28470 -42948 -28370 -42038
rect -27640 -42948 -27540 -42038
rect -26348 -42948 -26248 -41048
rect -24242 -42948 -24142 -41048
rect -22136 -42948 -22036 -41048
rect -20030 -42948 -19930 -41048
rect -17924 -42948 -17824 -41048
rect -15818 -42948 -15718 -41048
rect -13712 -42948 -13612 -41048
rect -11606 -42948 -11506 -41048
rect -9500 -42948 -9400 -41048
rect -7394 -42948 -7294 -41048
rect -5288 -42948 -5188 -41048
rect -3182 -42948 -3082 -41048
rect -1076 -42948 -976 -41048
rect 1030 -42948 1130 -41048
rect 3136 -42948 3236 -41048
rect 5242 -42948 5342 -41048
rect 7368 -41942 7468 -41048
rect 8160 -41942 8260 -41048
rect 7330 -42042 8260 -41942
rect 7368 -42948 7468 -42042
rect 8160 -42948 8260 -42042
rect -28470 -43048 8260 -42948
rect 26980 -42937 27052 -42936
rect 26980 -43001 26981 -42937
rect 27051 -43001 27052 -42937
rect 26980 -43002 27052 -43001
rect -28470 -43938 -28370 -43048
rect -27640 -43938 -27540 -43048
rect -28470 -44038 -27540 -43938
rect -28470 -44942 -28370 -44038
rect -27640 -44942 -27540 -44038
rect -26348 -44942 -26248 -43048
rect -24242 -44942 -24142 -43048
rect -22136 -44942 -22036 -43048
rect -20030 -44942 -19930 -43048
rect -17924 -44942 -17824 -43048
rect -15818 -44942 -15718 -43048
rect -13712 -44942 -13612 -43048
rect -11606 -44942 -11506 -43048
rect -9500 -44942 -9400 -43048
rect -28470 -45042 -9400 -44942
rect -8684 -44864 -8584 -44560
rect -8684 -44964 -8182 -44864
rect -7394 -44948 -7294 -43048
rect -5288 -44948 -5188 -43048
rect -3182 -44948 -3082 -43048
rect -1076 -44948 -976 -43048
rect 1030 -44948 1130 -43048
rect 3136 -44948 3236 -43048
rect 5242 -44948 5342 -43048
rect 7368 -43942 7468 -43048
rect 8160 -43942 8260 -43048
rect 7330 -44042 8260 -43942
rect 51344 -43984 53126 -43184
rect 7368 -44948 7468 -44042
rect 8160 -44948 8260 -44042
rect -28470 -45938 -28370 -45042
rect -27640 -45938 -27540 -45042
rect -28470 -46038 -27540 -45938
rect -28470 -46950 -28370 -46038
rect -27640 -46950 -27540 -46038
rect -26348 -46950 -26248 -45042
rect -24242 -46950 -24142 -45042
rect -22136 -46950 -22036 -45042
rect -20030 -46950 -19930 -45042
rect -17924 -46950 -17824 -45042
rect -15818 -46950 -15718 -45042
rect -13712 -46950 -13612 -45042
rect -11606 -46950 -11506 -45042
rect -28470 -47050 -11506 -46950
rect -10794 -46922 -10694 -46420
rect -10794 -47022 -10292 -46922
rect -28470 -47938 -28370 -47050
rect -27640 -47938 -27540 -47050
rect -28470 -48038 -27540 -47938
rect -28470 -48952 -28370 -48038
rect -27640 -48952 -27540 -48038
rect -26348 -48952 -26248 -47050
rect -24242 -48952 -24142 -47050
rect -22136 -48952 -22036 -47050
rect -20030 -48952 -19930 -47050
rect -17924 -48952 -17824 -47050
rect -15818 -48952 -15718 -47050
rect -28470 -49052 -15718 -48952
rect -15000 -48900 -14900 -48486
rect -15000 -49000 -14652 -48900
rect -28470 -49938 -28370 -49052
rect -27640 -49938 -27540 -49052
rect -28470 -50038 -27540 -49938
rect -28470 -50966 -28370 -50038
rect -27640 -50966 -27540 -50038
rect -26348 -50966 -26248 -49052
rect -24242 -50966 -24142 -49052
rect -22136 -50966 -22036 -49052
rect -20030 -50966 -19930 -49052
rect -17924 -50966 -17824 -49052
rect -15818 -50966 -15718 -49052
rect -28470 -51066 -15718 -50966
rect -28470 -51938 -28370 -51066
rect -27640 -51938 -27540 -51066
rect -28470 -52038 -27540 -51938
rect -28470 -52962 -28370 -52038
rect -27640 -52962 -27540 -52038
rect -26348 -52962 -26248 -51066
rect -24242 -52962 -24142 -51066
rect -22136 -52962 -22036 -51066
rect -20030 -52962 -19930 -51066
rect -17924 -52962 -17824 -51066
rect -28470 -53062 -17824 -52962
rect -28470 -53938 -28370 -53062
rect -27640 -53938 -27540 -53062
rect -28470 -54038 -27540 -53938
rect -28470 -54956 -28370 -54038
rect -27640 -54956 -27540 -54038
rect -26348 -54956 -26248 -53062
rect -24242 -54956 -24142 -53062
rect -22136 -54956 -22036 -53062
rect -20030 -54956 -19930 -53062
rect -28470 -55056 -19930 -54956
rect -19212 -54926 -19112 -54450
rect -19212 -55026 -18864 -54926
rect -28470 -55938 -28370 -55056
rect -27640 -55938 -27540 -55056
rect -28470 -56038 -27540 -55938
rect -28470 -56966 -28370 -56038
rect -27640 -56966 -27540 -56038
rect -26348 -56966 -26248 -55056
rect -24242 -56966 -24142 -55056
rect -22136 -56966 -22036 -55056
rect -20030 -56966 -19930 -55056
rect -28470 -57066 -19930 -56966
rect -28470 -57938 -28370 -57066
rect -27640 -57938 -27540 -57066
rect -28470 -58038 -27540 -57938
rect -28470 -58934 -28370 -58038
rect -27640 -58934 -27540 -58038
rect -26348 -58934 -26248 -57066
rect -24242 -58934 -24142 -57066
rect -22136 -58934 -22036 -57066
rect -20030 -58934 -19930 -57066
rect -28470 -59034 -19930 -58934
rect -28470 -59938 -28370 -59034
rect -27640 -59938 -27540 -59034
rect -28470 -60038 -27540 -59938
rect -28470 -60942 -28370 -60038
rect -27640 -60942 -27540 -60038
rect -26348 -60942 -26248 -59034
rect -24242 -60942 -24142 -59034
rect -22136 -60942 -22036 -59034
rect -20030 -60942 -19930 -59034
rect -28470 -61042 -19930 -60942
rect -28470 -61936 -28370 -61042
rect -27640 -61936 -27540 -61042
rect -26348 -61936 -26248 -61042
rect -24242 -61930 -24142 -61042
rect -22136 -61908 -22036 -61042
rect -20030 -61908 -19930 -61042
rect -24242 -61936 -23350 -61930
rect -22136 -61936 -21244 -61930
rect -20030 -61936 -19138 -61930
rect -28470 -62030 -19138 -61936
rect -28470 -62036 -19570 -62030
rect -18964 -63015 -18864 -55026
rect -17924 -61908 -17824 -53062
rect -17114 -52968 -17014 -52416
rect -17114 -53068 -16748 -52968
rect -17924 -62030 -17032 -61930
rect -18964 -63113 -18963 -63015
rect -18865 -63113 -18864 -63015
rect -16848 -63011 -16748 -53068
rect -15818 -61908 -15718 -51066
rect -15818 -62030 -14926 -61930
rect -16848 -63109 -16847 -63011
rect -16749 -63109 -16748 -63011
rect -14752 -63009 -14652 -49000
rect -13712 -61908 -13612 -47050
rect -12906 -48898 -12806 -48394
rect -12906 -48998 -12528 -48898
rect -13712 -62030 -12820 -61930
rect -14752 -63107 -14751 -63009
rect -14653 -63107 -14652 -63009
rect -14752 -63108 -14652 -63107
rect -12628 -63019 -12528 -48998
rect -11606 -61908 -11506 -47050
rect -10794 -48956 -10694 -48326
rect -10794 -49056 -10492 -48956
rect -11606 -62030 -10714 -61930
rect -16848 -63110 -16748 -63109
rect -18964 -63114 -18864 -63113
rect -12628 -63117 -12627 -63019
rect -12529 -63117 -12528 -63019
rect -10592 -63011 -10492 -49056
rect -10592 -63109 -10591 -63011
rect -10493 -63109 -10492 -63011
rect -10392 -63000 -10292 -47022
rect -9500 -61908 -9400 -45042
rect -8688 -47012 -8588 -46382
rect -8688 -47112 -8396 -47012
rect -9500 -62030 -8608 -61930
rect -10392 -63001 -9838 -63000
rect -10392 -63099 -9937 -63001
rect -9839 -63099 -9838 -63001
rect -10392 -63100 -9838 -63099
rect -8496 -63019 -8396 -47112
rect -10592 -63110 -10492 -63109
rect -12628 -63118 -12528 -63117
rect -8496 -63117 -8495 -63019
rect -8397 -63117 -8396 -63019
rect -8496 -63118 -8396 -63117
rect -8282 -63022 -8182 -44964
rect -7408 -45048 8260 -44948
rect -7394 -46948 -7294 -45048
rect -5288 -46948 -5188 -45048
rect -3182 -46948 -3082 -45048
rect -1076 -46948 -976 -45048
rect 1030 -46948 1130 -45048
rect 3136 -46948 3236 -45048
rect 5242 -46948 5342 -45048
rect 7368 -45942 7468 -45048
rect 8160 -45942 8260 -45048
rect 7330 -46042 8260 -45942
rect 7368 -46948 7468 -46042
rect 8160 -46948 8260 -46042
rect -7394 -47048 8260 -46948
rect -7394 -48948 -7294 -47048
rect -5288 -48948 -5188 -47048
rect -3182 -48948 -3082 -47048
rect -1076 -48948 -976 -47048
rect 1030 -48948 1130 -47048
rect 3136 -48948 3236 -47048
rect 5242 -48948 5342 -47048
rect 7368 -47942 7468 -47048
rect 8160 -47942 8260 -47048
rect 7330 -48042 8260 -47942
rect 7368 -48948 7468 -48042
rect 8160 -48948 8260 -48042
rect -7394 -49048 8260 -48948
rect -7394 -61908 -7294 -49048
rect -5288 -50948 -5188 -49048
rect -3182 -50948 -3082 -49048
rect -1076 -50948 -976 -49048
rect 1030 -50948 1130 -49048
rect 3136 -50948 3236 -49048
rect 5242 -50948 5342 -49048
rect 7368 -49942 7468 -49048
rect 8160 -49942 8260 -49048
rect 7330 -50042 8260 -49942
rect 7368 -50948 7468 -50042
rect 8160 -50948 8260 -50042
rect -5288 -51048 8260 -50948
rect -5288 -52948 -5188 -51048
rect -3182 -52948 -3082 -51048
rect -1076 -52948 -976 -51048
rect 1030 -52948 1130 -51048
rect 3136 -52948 3236 -51048
rect 5242 -52948 5342 -51048
rect 7368 -51942 7468 -51048
rect 8160 -51942 8260 -51048
rect 7330 -52042 8260 -51942
rect 7368 -52948 7468 -52042
rect 8160 -52948 8260 -52042
rect -5288 -52949 8264 -52948
rect -5288 -53047 8165 -52949
rect 8263 -53047 8264 -52949
rect -5288 -53048 8264 -53047
rect -5288 -54948 -5188 -53048
rect -3182 -54948 -3082 -53048
rect -1076 -54948 -976 -53048
rect 1030 -54948 1130 -53048
rect 3136 -54948 3236 -53048
rect 5242 -54948 5342 -53048
rect 7368 -53942 7468 -53048
rect 8160 -53942 8260 -53048
rect 7330 -54042 8260 -53942
rect 7368 -54948 7468 -54042
rect 8160 -54948 8260 -54042
rect -5288 -54949 8262 -54948
rect -5288 -55047 8163 -54949
rect 8261 -55047 8262 -54949
rect -5288 -55048 8262 -55047
rect -5288 -56948 -5188 -55048
rect -3182 -56948 -3082 -55048
rect -1076 -56948 -976 -55048
rect 1030 -56948 1130 -55048
rect 3136 -56948 3236 -55048
rect 5242 -56948 5342 -55048
rect 7368 -55942 7468 -55048
rect 8160 -55942 8260 -55048
rect 7330 -56042 8260 -55942
rect 7368 -56948 7468 -56042
rect 8160 -56948 8260 -56042
rect -5288 -57048 8260 -56948
rect -5288 -58948 -5188 -57048
rect -3182 -58948 -3082 -57048
rect -1076 -58948 -976 -57048
rect 1030 -58948 1130 -57048
rect 3136 -58948 3236 -57048
rect 5242 -58948 5342 -57048
rect 7368 -57942 7468 -57048
rect 8160 -57942 8260 -57048
rect 7330 -58042 8260 -57942
rect 7368 -58948 7468 -58042
rect 8160 -58948 8260 -58042
rect -5288 -59048 8260 -58948
rect -5288 -60968 -5188 -59048
rect -3182 -60968 -3082 -59048
rect -1076 -60968 -976 -59048
rect 1030 -60968 1130 -59048
rect 3136 -60968 3236 -59048
rect 5242 -60968 5342 -59048
rect 7368 -59942 7468 -59048
rect 8160 -59942 8260 -59048
rect 49716 -58404 51344 -58380
rect 49716 -59156 50568 -58404
rect 51320 -59156 51344 -58404
rect 49716 -59180 51344 -59156
rect 7330 -60042 8260 -59942
rect 7368 -60968 7468 -60042
rect 8160 -60968 8260 -60042
rect -5288 -61068 8260 -60968
rect -5288 -61908 -5188 -61068
rect -3182 -61908 -3082 -61068
rect -1076 -61908 -976 -61068
rect 1030 -61908 1130 -61068
rect 3136 -61908 3236 -61068
rect 5242 -61930 5342 -61068
rect 7368 -61930 7468 -61068
rect -7394 -62030 -6502 -61930
rect -5288 -61936 7476 -61930
rect 8160 -61936 8260 -61068
rect -5288 -62030 8260 -61936
rect 5202 -62036 8260 -62030
rect 8160 -62122 8260 -62036
rect -8282 -63023 -7828 -63022
rect -8282 -63121 -7927 -63023
rect -7829 -63121 -7828 -63023
rect -8282 -63122 -7828 -63121
rect -27764 -65036 7040 -64348
rect 7728 -65036 8854 -64348
rect -26889 -69716 -26223 -69222
rect -22859 -69716 -22193 -69222
rect -18837 -69716 -18171 -69222
rect -14853 -69716 -14187 -69222
rect -10909 -69716 -10243 -69222
rect -6853 -69716 -6187 -69222
rect -2875 -69716 -2209 -69222
rect 1153 -69716 1819 -69222
rect 5131 -69716 5797 -69222
rect 9356 -69716 11076 -69714
rect -27762 -69738 11076 -69716
rect -27762 -70490 10300 -69738
rect 11052 -70490 11076 -69738
rect -27762 -70514 11076 -70490
rect -27762 -70516 10276 -70514
rect -26889 -70941 -26223 -70516
rect -22859 -70875 -22193 -70516
rect -18837 -70901 -18171 -70516
rect -14853 -70913 -14187 -70516
rect -10909 -70853 -10243 -70516
rect -6853 -70859 -6187 -70516
rect -2875 -70877 -2209 -70516
rect 1153 -70889 1819 -70516
rect 5131 -70871 5797 -70516
rect -27760 -75178 7728 -75160
rect -27760 -75818 7064 -75178
rect 7704 -75818 7728 -75178
rect -27760 -75848 7728 -75818
<< via4 >>
rect 8788 -28378 9588 -27578
rect 50552 -28378 51352 -27578
rect 50576 -39456 51328 -38704
rect 50544 -43984 51344 -43184
rect 9250 -56724 9554 -56598
rect 9250 -57518 9372 -56724
rect 9372 -57518 9436 -56724
rect 9436 -57518 9554 -56724
rect 9250 -57594 9554 -57518
rect 10276 -58408 11076 -58378
rect 10276 -58514 10294 -58408
rect 10294 -58514 11076 -58408
rect 10276 -59178 11076 -58514
rect 50568 -59156 51320 -58404
rect 7040 -65036 7728 -64348
rect 8854 -65036 9542 -64348
rect 10300 -70490 11052 -69738
rect 7064 -75818 7704 -75178
<< metal5 >>
rect 8764 -27578 9612 -27554
rect 8764 -28378 8788 -27578
rect 9588 -28378 9612 -27578
rect 8764 -28402 9612 -28378
rect 50528 -27578 51376 -27554
rect 50528 -28378 50552 -27578
rect 51352 -28378 51376 -27578
rect 50528 -28402 51376 -28378
rect 8788 -56598 9588 -28402
rect 50552 -38704 51352 -28402
rect 50552 -39456 50576 -38704
rect 51328 -39456 51352 -38704
rect 50552 -39480 51352 -39456
rect 50520 -43184 51368 -43160
rect 50520 -43984 50544 -43184
rect 51344 -43984 51368 -43184
rect 50520 -44008 51368 -43984
rect 8788 -57594 9250 -56598
rect 9554 -57594 9588 -56598
rect 7016 -64348 7752 -64324
rect 7016 -65036 7040 -64348
rect 7728 -65036 7752 -64348
rect 7016 -65060 7752 -65036
rect 8788 -64348 9588 -57594
rect 10252 -58378 11100 -58354
rect 10252 -59178 10276 -58378
rect 11076 -59178 11100 -58378
rect 10252 -59202 11100 -59178
rect 50544 -58404 51344 -44008
rect 50544 -59156 50568 -58404
rect 51320 -59156 51344 -58404
rect 50544 -59180 51344 -59156
rect 8788 -65036 8854 -64348
rect 9542 -65036 9588 -64348
rect 7040 -75178 7728 -65060
rect 8788 -65088 9588 -65036
rect 10276 -69738 11076 -59202
rect 10276 -70490 10300 -69738
rect 11052 -70490 11076 -69738
rect 10276 -70514 11076 -70490
rect 7040 -75818 7064 -75178
rect 7704 -75818 7728 -75178
rect 7040 -75842 7728 -75818
use amux_2to1  amux_2to1_17 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/amux_2to1
timestamp 1624127230
transform 1 0 -28122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_16
timestamp 1624127230
transform 1 0 -24122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_15
timestamp 1624127230
transform 1 0 -20122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_14
timestamp 1624127230
transform 1 0 -16122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_13
timestamp 1624127230
transform 1 0 -12122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_12
timestamp 1624127230
transform 1 0 -8122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_11
timestamp 1624127230
transform 1 0 -4122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_10
timestamp 1624127230
transform 1 0 -122 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_9
timestamp 1624127230
transform 1 0 3878 0 -1 -72108
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_0
timestamp 1624127230
transform 1 0 -28122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_1
timestamp 1624127230
transform 1 0 -24122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_2
timestamp 1624127230
transform 1 0 -20122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_3
timestamp 1624127230
transform 1 0 -16122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_4
timestamp 1624127230
transform 1 0 -12122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_5
timestamp 1624127230
transform 1 0 -8122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_6
timestamp 1624127230
transform 1 0 -4122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_7
timestamp 1624127230
transform 1 0 -122 0 1 -68088
box -114 -1800 2840 3740
use amux_2to1  amux_2to1_8
timestamp 1624127230
transform 1 0 3878 0 1 -68088
box -114 -1800 2840 3740
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_17
timestamp 1624127230
transform 1 0 -28385 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_16
timestamp 1624127230
transform 1 0 -28385 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_18
timestamp 1624127230
transform 1 0 -26279 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_19
timestamp 1624127230
transform 1 0 -26279 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_36
timestamp 1624127230
transform 1 0 -24173 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_37
timestamp 1624127230
transform 1 0 -24173 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_54
timestamp 1624127230
transform 1 0 -22067 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_55
timestamp 1624127230
transform 1 0 -22067 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_73
timestamp 1624127230
transform 1 0 -19961 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_72
timestamp 1624127230
transform 1 0 -19961 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_91
timestamp 1624127230
transform 1 0 -17855 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_90
timestamp 1624127230
transform 1 0 -17855 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_109
timestamp 1624127230
transform 1 0 -15749 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_108
timestamp 1624127230
transform 1 0 -15749 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_127
timestamp 1624127230
transform 1 0 -13643 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_126
timestamp 1624127230
transform 1 0 -13643 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_145
timestamp 1624127230
transform 1 0 -11537 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_144
timestamp 1624127230
transform 1 0 -11537 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_163
timestamp 1624127230
transform 1 0 -9431 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_162
timestamp 1624127230
transform 1 0 -9431 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_181
timestamp 1624127230
transform 1 0 -7325 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_180
timestamp 1624127230
transform 1 0 -7325 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_199
timestamp 1624127230
transform 1 0 -5219 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_198
timestamp 1624127230
transform 1 0 -5219 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_217
timestamp 1624127230
transform 1 0 -3113 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_216
timestamp 1624127230
transform 1 0 -3113 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_235
timestamp 1624127230
transform 1 0 -1007 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_234
timestamp 1624127230
transform 1 0 -1007 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_253
timestamp 1624127230
transform 1 0 1099 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_252
timestamp 1624127230
transform 1 0 1099 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_271
timestamp 1624127230
transform 1 0 3205 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_270
timestamp 1624127230
transform 1 0 3205 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_289
timestamp 1624127230
transform 1 0 5311 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_288
timestamp 1624127230
transform 1 0 5311 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_307
timestamp 1624127230
transform 1 0 7417 0 1 -60006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_306
timestamp 1624127230
transform 1 0 7417 0 1 -62006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_15
timestamp 1624127230
transform 1 0 -28385 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_20
timestamp 1624127230
transform 1 0 -26279 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_14
timestamp 1624127230
transform 1 0 -28385 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_21
timestamp 1624127230
transform 1 0 -26279 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_13
timestamp 1624127230
transform 1 0 -28385 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_22
timestamp 1624127230
transform 1 0 -26279 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_38
timestamp 1624127230
transform 1 0 -24173 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_39
timestamp 1624127230
transform 1 0 -24173 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_40
timestamp 1624127230
transform 1 0 -24173 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_56
timestamp 1624127230
transform 1 0 -22067 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_57
timestamp 1624127230
transform 1 0 -22067 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_58
timestamp 1624127230
transform 1 0 -22067 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_74
timestamp 1624127230
transform 1 0 -19961 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_75
timestamp 1624127230
transform 1 0 -19961 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_76
timestamp 1624127230
transform 1 0 -19961 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_92
timestamp 1624127230
transform 1 0 -17855 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_93
timestamp 1624127230
transform 1 0 -17855 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_94
timestamp 1624127230
transform 1 0 -17855 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_110
timestamp 1624127230
transform 1 0 -15749 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_128
timestamp 1624127230
transform 1 0 -13643 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_111
timestamp 1624127230
transform 1 0 -15749 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_129
timestamp 1624127230
transform 1 0 -13643 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_112
timestamp 1624127230
transform 1 0 -15749 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_130
timestamp 1624127230
transform 1 0 -13643 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_146
timestamp 1624127230
transform 1 0 -11537 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_147
timestamp 1624127230
transform 1 0 -11537 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_148
timestamp 1624127230
transform 1 0 -11537 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_164
timestamp 1624127230
transform 1 0 -9431 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_165
timestamp 1624127230
transform 1 0 -9431 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_166
timestamp 1624127230
transform 1 0 -9431 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_182
timestamp 1624127230
transform 1 0 -7325 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_183
timestamp 1624127230
transform 1 0 -7325 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_184
timestamp 1624127230
transform 1 0 -7325 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_200
timestamp 1624127230
transform 1 0 -5219 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_201
timestamp 1624127230
transform 1 0 -5219 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_202
timestamp 1624127230
transform 1 0 -5219 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_218
timestamp 1624127230
transform 1 0 -3113 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_219
timestamp 1624127230
transform 1 0 -3113 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_220
timestamp 1624127230
transform 1 0 -3113 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_236
timestamp 1624127230
transform 1 0 -1007 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_254
timestamp 1624127230
transform 1 0 1099 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_237
timestamp 1624127230
transform 1 0 -1007 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_255
timestamp 1624127230
transform 1 0 1099 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_238
timestamp 1624127230
transform 1 0 -1007 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_256
timestamp 1624127230
transform 1 0 1099 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_272
timestamp 1624127230
transform 1 0 3205 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_273
timestamp 1624127230
transform 1 0 3205 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_274
timestamp 1624127230
transform 1 0 3205 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_290
timestamp 1624127230
transform 1 0 5311 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_291
timestamp 1624127230
transform 1 0 5311 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_292
timestamp 1624127230
transform 1 0 5311 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_308
timestamp 1624127230
transform 1 0 7417 0 1 -58006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_309
timestamp 1624127230
transform 1 0 7417 0 1 -56006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_310
timestamp 1624127230
transform 1 0 7417 0 1 -54006
box -850 -800 849 800
use sky130_fd_pr__pfet_01v8_hvt_SCHXZ7  sky130_fd_pr__pfet_01v8_hvt_SCHXZ7_0
timestamp 1624127230
transform 1 0 11201 0 1 -57122
box -941 -419 941 419
use sky130_fd_pr__nfet_01v8_N6QVV6  sky130_fd_pr__nfet_01v8_N6QVV6_0
timestamp 1624127230
transform 1 0 11201 0 1 -57946
box -941 -310 941 310
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_12
timestamp 1624127230
transform 1 0 -28385 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_23
timestamp 1624127230
transform 1 0 -26279 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_41
timestamp 1624127230
transform 1 0 -24173 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_59
timestamp 1624127230
transform 1 0 -22067 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_77
timestamp 1624127230
transform 1 0 -19961 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_95
timestamp 1624127230
transform 1 0 -17855 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_113
timestamp 1624127230
transform 1 0 -15749 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_131
timestamp 1624127230
transform 1 0 -13643 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_149
timestamp 1624127230
transform 1 0 -11537 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_167
timestamp 1624127230
transform 1 0 -9431 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_185
timestamp 1624127230
transform 1 0 -7325 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_203
timestamp 1624127230
transform 1 0 -5219 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_221
timestamp 1624127230
transform 1 0 -3113 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_239
timestamp 1624127230
transform 1 0 -1007 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_257
timestamp 1624127230
transform 1 0 1099 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_275
timestamp 1624127230
transform 1 0 3205 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_293
timestamp 1624127230
transform 1 0 5311 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_311
timestamp 1624127230
transform 1 0 7417 0 1 -52006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_11
timestamp 1624127230
transform 1 0 -28385 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_24
timestamp 1624127230
transform 1 0 -26279 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_42
timestamp 1624127230
transform 1 0 -24173 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_60
timestamp 1624127230
transform 1 0 -22067 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_78
timestamp 1624127230
transform 1 0 -19961 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_96
timestamp 1624127230
transform 1 0 -17855 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_114
timestamp 1624127230
transform 1 0 -15749 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_132
timestamp 1624127230
transform 1 0 -13643 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_150
timestamp 1624127230
transform 1 0 -11537 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_168
timestamp 1624127230
transform 1 0 -9431 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_186
timestamp 1624127230
transform 1 0 -7325 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_204
timestamp 1624127230
transform 1 0 -5219 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_222
timestamp 1624127230
transform 1 0 -3113 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_240
timestamp 1624127230
transform 1 0 -1007 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_258
timestamp 1624127230
transform 1 0 1099 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_276
timestamp 1624127230
transform 1 0 3205 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_294
timestamp 1624127230
transform 1 0 5311 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_312
timestamp 1624127230
transform 1 0 7417 0 1 -50006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_10
timestamp 1624127230
transform 1 0 -28385 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_25
timestamp 1624127230
transform 1 0 -26279 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_43
timestamp 1624127230
transform 1 0 -24173 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_61
timestamp 1624127230
transform 1 0 -22067 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_79
timestamp 1624127230
transform 1 0 -19961 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_97
timestamp 1624127230
transform 1 0 -17855 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_115
timestamp 1624127230
transform 1 0 -15749 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_133
timestamp 1624127230
transform 1 0 -13643 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_151
timestamp 1624127230
transform 1 0 -11537 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_169
timestamp 1624127230
transform 1 0 -9431 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_187
timestamp 1624127230
transform 1 0 -7325 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_205
timestamp 1624127230
transform 1 0 -5219 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_223
timestamp 1624127230
transform 1 0 -3113 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_241
timestamp 1624127230
transform 1 0 -1007 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_259
timestamp 1624127230
transform 1 0 1099 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_277
timestamp 1624127230
transform 1 0 3205 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_295
timestamp 1624127230
transform 1 0 5311 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_313
timestamp 1624127230
transform 1 0 7417 0 1 -48006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_9
timestamp 1624127230
transform 1 0 -28385 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_26
timestamp 1624127230
transform 1 0 -26279 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_44
timestamp 1624127230
transform 1 0 -24173 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_62
timestamp 1624127230
transform 1 0 -22067 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_80
timestamp 1624127230
transform 1 0 -19961 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_98
timestamp 1624127230
transform 1 0 -17855 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_116
timestamp 1624127230
transform 1 0 -15749 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_134
timestamp 1624127230
transform 1 0 -13643 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_152
timestamp 1624127230
transform 1 0 -11537 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_170
timestamp 1624127230
transform 1 0 -9431 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_188
timestamp 1624127230
transform 1 0 -7325 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_206
timestamp 1624127230
transform 1 0 -5219 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_224
timestamp 1624127230
transform 1 0 -3113 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_242
timestamp 1624127230
transform 1 0 -1007 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_260
timestamp 1624127230
transform 1 0 1099 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_278
timestamp 1624127230
transform 1 0 3205 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_296
timestamp 1624127230
transform 1 0 5311 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_314
timestamp 1624127230
transform 1 0 7417 0 1 -46006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_8
timestamp 1624127230
transform 1 0 -28385 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_27
timestamp 1624127230
transform 1 0 -26279 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_45
timestamp 1624127230
transform 1 0 -24173 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_63
timestamp 1624127230
transform 1 0 -22067 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_81
timestamp 1624127230
transform 1 0 -19961 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_99
timestamp 1624127230
transform 1 0 -17855 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_117
timestamp 1624127230
transform 1 0 -15749 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_135
timestamp 1624127230
transform 1 0 -13643 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_153
timestamp 1624127230
transform 1 0 -11537 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_171
timestamp 1624127230
transform 1 0 -9431 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_189
timestamp 1624127230
transform 1 0 -7325 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_207
timestamp 1624127230
transform 1 0 -5219 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_225
timestamp 1624127230
transform 1 0 -3113 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_243
timestamp 1624127230
transform 1 0 -1007 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_261
timestamp 1624127230
transform 1 0 1099 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_279
timestamp 1624127230
transform 1 0 3205 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_297
timestamp 1624127230
transform 1 0 5311 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_315
timestamp 1624127230
transform 1 0 7417 0 1 -44006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_7
timestamp 1624127230
transform 1 0 -28385 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_28
timestamp 1624127230
transform 1 0 -26279 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_46
timestamp 1624127230
transform 1 0 -24173 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_64
timestamp 1624127230
transform 1 0 -22067 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_82
timestamp 1624127230
transform 1 0 -19961 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_100
timestamp 1624127230
transform 1 0 -17855 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_118
timestamp 1624127230
transform 1 0 -15749 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_136
timestamp 1624127230
transform 1 0 -13643 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_154
timestamp 1624127230
transform 1 0 -11537 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_172
timestamp 1624127230
transform 1 0 -9431 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_190
timestamp 1624127230
transform 1 0 -7325 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_208
timestamp 1624127230
transform 1 0 -5219 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_226
timestamp 1624127230
transform 1 0 -3113 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_244
timestamp 1624127230
transform 1 0 -1007 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_262
timestamp 1624127230
transform 1 0 1099 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_280
timestamp 1624127230
transform 1 0 3205 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_298
timestamp 1624127230
transform 1 0 5311 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_316
timestamp 1624127230
transform 1 0 7417 0 1 -42006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_6
timestamp 1624127230
transform 1 0 -28385 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_29
timestamp 1624127230
transform 1 0 -26279 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_5
timestamp 1624127230
transform 1 0 -28385 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_30
timestamp 1624127230
transform 1 0 -26279 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_47
timestamp 1624127230
transform 1 0 -24173 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_48
timestamp 1624127230
transform 1 0 -24173 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_65
timestamp 1624127230
transform 1 0 -22067 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_66
timestamp 1624127230
transform 1 0 -22067 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_83
timestamp 1624127230
transform 1 0 -19961 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_84
timestamp 1624127230
transform 1 0 -19961 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_101
timestamp 1624127230
transform 1 0 -17855 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_102
timestamp 1624127230
transform 1 0 -17855 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_119
timestamp 1624127230
transform 1 0 -15749 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_120
timestamp 1624127230
transform 1 0 -15749 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_137
timestamp 1624127230
transform 1 0 -13643 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_138
timestamp 1624127230
transform 1 0 -13643 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_155
timestamp 1624127230
transform 1 0 -11537 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_156
timestamp 1624127230
transform 1 0 -11537 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_173
timestamp 1624127230
transform 1 0 -9431 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_174
timestamp 1624127230
transform 1 0 -9431 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_191
timestamp 1624127230
transform 1 0 -7325 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_192
timestamp 1624127230
transform 1 0 -7325 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_209
timestamp 1624127230
transform 1 0 -5219 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_210
timestamp 1624127230
transform 1 0 -5219 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_227
timestamp 1624127230
transform 1 0 -3113 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_228
timestamp 1624127230
transform 1 0 -3113 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_245
timestamp 1624127230
transform 1 0 -1007 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_246
timestamp 1624127230
transform 1 0 -1007 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_263
timestamp 1624127230
transform 1 0 1099 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_264
timestamp 1624127230
transform 1 0 1099 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_281
timestamp 1624127230
transform 1 0 3205 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_282
timestamp 1624127230
transform 1 0 3205 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_299
timestamp 1624127230
transform 1 0 5311 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_300
timestamp 1624127230
transform 1 0 5311 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_317
timestamp 1624127230
transform 1 0 7417 0 1 -40006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_318
timestamp 1624127230
transform 1 0 7417 0 1 -38006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_4
timestamp 1624127230
transform 1 0 -28385 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_31
timestamp 1624127230
transform 1 0 -26279 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_49
timestamp 1624127230
transform 1 0 -24173 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_67
timestamp 1624127230
transform 1 0 -22067 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_85
timestamp 1624127230
transform 1 0 -19961 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_103
timestamp 1624127230
transform 1 0 -17855 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_121
timestamp 1624127230
transform 1 0 -15749 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_139
timestamp 1624127230
transform 1 0 -13643 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_157
timestamp 1624127230
transform 1 0 -11537 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_175
timestamp 1624127230
transform 1 0 -9431 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_193
timestamp 1624127230
transform 1 0 -7325 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_211
timestamp 1624127230
transform 1 0 -5219 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_229
timestamp 1624127230
transform 1 0 -3113 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_247
timestamp 1624127230
transform 1 0 -1007 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_265
timestamp 1624127230
transform 1 0 1099 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_283
timestamp 1624127230
transform 1 0 3205 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_301
timestamp 1624127230
transform 1 0 5311 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_319
timestamp 1624127230
transform 1 0 7417 0 1 -36006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_3
timestamp 1624127230
transform 1 0 -28385 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_32
timestamp 1624127230
transform 1 0 -26279 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_50
timestamp 1624127230
transform 1 0 -24173 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_68
timestamp 1624127230
transform 1 0 -22067 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_86
timestamp 1624127230
transform 1 0 -19961 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_104
timestamp 1624127230
transform 1 0 -17855 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_122
timestamp 1624127230
transform 1 0 -15749 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_140
timestamp 1624127230
transform 1 0 -13643 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_158
timestamp 1624127230
transform 1 0 -11537 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_176
timestamp 1624127230
transform 1 0 -9431 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_194
timestamp 1624127230
transform 1 0 -7325 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_212
timestamp 1624127230
transform 1 0 -5219 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_230
timestamp 1624127230
transform 1 0 -3113 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_248
timestamp 1624127230
transform 1 0 -1007 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_266
timestamp 1624127230
transform 1 0 1099 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_284
timestamp 1624127230
transform 1 0 3205 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_302
timestamp 1624127230
transform 1 0 5311 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_320
timestamp 1624127230
transform 1 0 7417 0 1 -34006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_2
timestamp 1624127230
transform 1 0 -28385 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_33
timestamp 1624127230
transform 1 0 -26279 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_51
timestamp 1624127230
transform 1 0 -24173 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_69
timestamp 1624127230
transform 1 0 -22067 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_87
timestamp 1624127230
transform 1 0 -19961 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_105
timestamp 1624127230
transform 1 0 -17855 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_123
timestamp 1624127230
transform 1 0 -15749 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_141
timestamp 1624127230
transform 1 0 -13643 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_159
timestamp 1624127230
transform 1 0 -11537 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_177
timestamp 1624127230
transform 1 0 -9431 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_195
timestamp 1624127230
transform 1 0 -7325 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_213
timestamp 1624127230
transform 1 0 -5219 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_231
timestamp 1624127230
transform 1 0 -3113 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_249
timestamp 1624127230
transform 1 0 -1007 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_267
timestamp 1624127230
transform 1 0 1099 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_285
timestamp 1624127230
transform 1 0 3205 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_303
timestamp 1624127230
transform 1 0 5311 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_321
timestamp 1624127230
transform 1 0 7417 0 1 -32006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_1
timestamp 1624127230
transform 1 0 -28385 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_34
timestamp 1624127230
transform 1 0 -26279 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_52
timestamp 1624127230
transform 1 0 -24173 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_70
timestamp 1624127230
transform 1 0 -22067 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_88
timestamp 1624127230
transform 1 0 -19961 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_106
timestamp 1624127230
transform 1 0 -17855 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_124
timestamp 1624127230
transform 1 0 -15749 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_142
timestamp 1624127230
transform 1 0 -13643 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_160
timestamp 1624127230
transform 1 0 -11537 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_178
timestamp 1624127230
transform 1 0 -9431 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_196
timestamp 1624127230
transform 1 0 -7325 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_214
timestamp 1624127230
transform 1 0 -5219 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_232
timestamp 1624127230
transform 1 0 -3113 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_250
timestamp 1624127230
transform 1 0 -1007 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_268
timestamp 1624127230
transform 1 0 1099 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_286
timestamp 1624127230
transform 1 0 3205 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_304
timestamp 1624127230
transform 1 0 5311 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_322
timestamp 1624127230
transform 1 0 7417 0 1 -30006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_0
timestamp 1624127230
transform 1 0 -28385 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_35
timestamp 1624127230
transform 1 0 -26279 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_53
timestamp 1624127230
transform 1 0 -24173 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_71
timestamp 1624127230
transform 1 0 -22067 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_89
timestamp 1624127230
transform 1 0 -19961 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_107
timestamp 1624127230
transform 1 0 -17855 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_125
timestamp 1624127230
transform 1 0 -15749 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_143
timestamp 1624127230
transform 1 0 -13643 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_161
timestamp 1624127230
transform 1 0 -11537 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_179
timestamp 1624127230
transform 1 0 -9431 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_197
timestamp 1624127230
transform 1 0 -7325 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_215
timestamp 1624127230
transform 1 0 -5219 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_233
timestamp 1624127230
transform 1 0 -3113 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_251
timestamp 1624127230
transform 1 0 -1007 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_269
timestamp 1624127230
transform 1 0 1099 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_287
timestamp 1624127230
transform 1 0 3205 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_305
timestamp 1624127230
transform 1 0 5311 0 1 -28006
box -850 -800 849 800
use sky130_fd_pr__cap_mim_m3_1_BZ3RER  sky130_fd_pr__cap_mim_m3_1_BZ3RER_323
timestamp 1624127230
transform 1 0 7417 0 1 -28006
box -850 -800 849 800
use se_fold_casc_wide_swing_ota  se_fold_casc_wide_swing_ota_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/se_fold_casc_wide_swing_ota
timestamp 1624132412
transform 1 0 25444 0 1 -31978
box -15168 -27258 25000 4400
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624127230
transform -1 0 12456 0 1 -57802
box -38 -48 314 592
use latched_comparator_folded  latched_comparator_folded_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/latched_comparator_folded
timestamp 1624127230
transform 1 0 55478 0 1 -40970
box -3400 -3014 3047 2278
<< labels >>
flabel metal3 -25220 -63116 -25188 -63092 1 FreeSans 480 0 0 0 c7m
flabel metal3 -18928 -63224 -18910 -63206 1 FreeSans 480 0 0 0 c6m
flabel metal3 -16804 -63244 -16796 -63228 1 FreeSans 480 0 0 0 c5m
flabel metal3 -14718 -63246 -14704 -63230 1 FreeSans 480 0 0 0 c4m
flabel metal3 -12590 -63222 -12576 -63208 1 FreeSans 480 0 0 0 c3m
flabel metal3 -8458 -63254 -8442 -63236 1 FreeSans 480 0 0 0 c1m
flabel metal3 -10548 -63244 -10520 -63220 1 FreeSans 480 0 0 0 c2m
flabel metal3 -9900 -63276 -9878 -63242 1 FreeSans 480 0 0 0 cdumm
flabel metal3 -7508 -63088 -7478 -63062 1 FreeSans 480 0 0 0 c0m
flabel metal4 -27544 -70138 -27514 -70094 1 FreeSans 480 0 0 0 VSS
flabel metal4 -27740 -64374 -27728 -64364 1 FreeSans 480 0 0 0 VDD
flabel metal3 -28160 -74900 -28146 -74892 1 FreeSans 480 0 0 0 vref
flabel metal3 -28452 -72922 -28438 -72906 1 FreeSans 480 0 0 0 vlow
flabel metal3 -28232 -67966 -28214 -67946 1 FreeSans 480 0 0 0 vin
flabel metal3 12544 -58056 12562 -58044 1 FreeSans 480 0 0 0 sample
flabel metal2 12200 -57048 12212 -57040 1 FreeSans 480 0 0 0 adc_run
flabel metal1 -28342 -72610 -28336 -72600 1 FreeSans 480 0 0 0 q7
flabel metal1 -24328 -72616 -24316 -72604 1 FreeSans 480 0 0 0 q6
flabel metal1 -20346 -72616 -20340 -72608 1 FreeSans 480 0 0 0 q5
flabel metal1 -16352 -72620 -16346 -72608 1 FreeSans 480 0 0 0 q4
flabel metal1 -12382 -72614 -12370 -72604 1 FreeSans 480 0 0 0 q3
flabel metal1 -8362 -72620 -8352 -72608 1 FreeSans 480 0 0 0 q2
flabel metal1 -356 -72608 -350 -72602 1 FreeSans 480 0 0 0 q1
flabel metal1 3634 -72616 3644 -72606 1 FreeSans 480 0 0 0 q0
flabel metal1 15262 -56936 15270 -56922 1 FreeSans 480 0 0 0 ibiasn
flabel metal3 10682 -52044 10722 -52028 1 FreeSans 480 0 0 0 vcom
flabel metal2 27012 -43058 27020 -43048 1 FreeSans 480 0 0 0 vcom_buf
flabel metal2 52036 -40050 52042 -40042 1 FreeSans 480 0 0 0 ibiasp
flabel metal2 52026 -42516 52034 -42508 1 FreeSans 480 0 0 0 adc_clk
flabel metal2 58410 -41968 58422 -41960 1 FreeSans 480 0 0 0 comp_out
flabel metal2 58400 -42168 58406 -42162 1 FreeSans 480 0 0 0 comp_outm
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< error_p >>
rect -1129 1100 -1089 1700
rect -1069 1100 -1029 1700
rect -410 1100 -370 1700
rect -350 1100 -310 1700
rect 309 1100 349 1700
rect 369 1100 409 1700
rect 1028 1100 1068 1700
rect 1088 1100 1128 1700
rect -1129 400 -1089 1000
rect -1069 400 -1029 1000
rect -410 400 -370 1000
rect -350 400 -310 1000
rect 309 400 349 1000
rect 369 400 409 1000
rect 1028 400 1068 1000
rect 1088 400 1128 1000
rect -1129 -300 -1089 300
rect -1069 -300 -1029 300
rect -410 -300 -370 300
rect -350 -300 -310 300
rect 309 -300 349 300
rect 369 -300 409 300
rect 1028 -300 1068 300
rect 1088 -300 1128 300
rect -1129 -1000 -1089 -400
rect -1069 -1000 -1029 -400
rect -410 -1000 -370 -400
rect -350 -1000 -310 -400
rect 309 -1000 349 -400
rect 369 -1000 409 -400
rect 1028 -1000 1068 -400
rect 1088 -1000 1128 -400
rect -1129 -1700 -1089 -1100
rect -1069 -1700 -1029 -1100
rect -410 -1700 -370 -1100
rect -350 -1700 -310 -1100
rect 309 -1700 349 -1100
rect 369 -1700 409 -1100
rect 1028 -1700 1068 -1100
rect 1088 -1700 1128 -1100
<< metal3 >>
rect -1788 1584 -1089 1700
rect -1788 1212 -1173 1584
rect -1109 1212 -1089 1584
rect -1788 1100 -1089 1212
rect -1069 1582 -370 1700
rect -1069 1212 -454 1582
rect -390 1212 -370 1582
rect -1069 1100 -370 1212
rect -350 1582 349 1700
rect -350 1212 265 1582
rect 329 1212 349 1582
rect -350 1100 349 1212
rect 369 1582 1068 1700
rect 369 1212 984 1582
rect 1048 1212 1068 1582
rect 369 1100 1068 1212
rect 1088 1582 1787 1700
rect 1088 1212 1703 1582
rect 1767 1212 1787 1582
rect 1088 1100 1787 1212
rect -1788 882 -1089 1000
rect -1788 514 -1173 882
rect -1109 514 -1089 882
rect -1788 400 -1089 514
rect -1069 882 -370 1000
rect -1069 514 -454 882
rect -390 514 -370 882
rect -1069 400 -370 514
rect -350 882 349 1000
rect -350 514 265 882
rect 329 514 349 882
rect -350 400 349 514
rect 369 882 1068 1000
rect 369 514 984 882
rect 1048 514 1068 882
rect 369 400 1068 514
rect 1088 882 1787 1000
rect 1088 514 1703 882
rect 1767 514 1787 882
rect 1088 400 1787 514
rect -1788 182 -1089 300
rect -1788 -186 -1173 182
rect -1109 -186 -1089 182
rect -1788 -300 -1089 -186
rect -1069 182 -370 300
rect -1069 -186 -454 182
rect -390 -186 -370 182
rect -1069 -300 -370 -186
rect -350 182 349 300
rect -350 -186 265 182
rect 329 -186 349 182
rect -350 -300 349 -186
rect 369 182 1068 300
rect 369 -186 984 182
rect 1048 -186 1068 182
rect 369 -300 1068 -186
rect 1088 182 1787 300
rect 1088 -186 1703 182
rect 1767 -186 1787 182
rect 1088 -300 1787 -186
rect -1788 -518 -1089 -400
rect -1788 -886 -1173 -518
rect -1109 -886 -1089 -518
rect -1788 -1000 -1089 -886
rect -1069 -518 -370 -400
rect -1069 -886 -454 -518
rect -390 -886 -370 -518
rect -1069 -1000 -370 -886
rect -350 -518 349 -400
rect -350 -886 265 -518
rect 329 -886 349 -518
rect -350 -1000 349 -886
rect 369 -518 1068 -400
rect 369 -886 984 -518
rect 1048 -886 1068 -518
rect 369 -1000 1068 -886
rect 1088 -518 1787 -400
rect 1088 -886 1703 -518
rect 1767 -886 1787 -518
rect 1088 -1000 1787 -886
rect -1788 -1218 -1089 -1100
rect -1788 -1586 -1173 -1218
rect -1109 -1586 -1089 -1218
rect -1788 -1700 -1089 -1586
rect -1069 -1218 -370 -1100
rect -1069 -1586 -454 -1218
rect -390 -1586 -370 -1218
rect -1069 -1700 -370 -1586
rect -350 -1218 349 -1100
rect -350 -1586 265 -1218
rect 329 -1586 349 -1218
rect -350 -1700 349 -1586
rect 369 -1218 1068 -1100
rect 369 -1586 984 -1218
rect 1048 -1586 1068 -1218
rect 369 -1700 1068 -1586
rect 1088 -1218 1787 -1100
rect 1088 -1586 1703 -1218
rect 1767 -1586 1787 -1218
rect 1088 -1700 1787 -1586
<< via3 >>
rect -1173 1212 -1109 1584
rect -454 1212 -390 1582
rect 265 1212 329 1582
rect 984 1212 1048 1582
rect 1703 1212 1767 1582
rect -1173 514 -1109 882
rect -454 514 -390 882
rect 265 514 329 882
rect 984 514 1048 882
rect 1703 514 1767 882
rect -1173 -186 -1109 182
rect -454 -186 -390 182
rect 265 -186 329 182
rect 984 -186 1048 182
rect 1703 -186 1767 182
rect -1173 -886 -1109 -518
rect -454 -886 -390 -518
rect 265 -886 329 -518
rect 984 -886 1048 -518
rect 1703 -886 1767 -518
rect -1173 -1586 -1109 -1218
rect -454 -1586 -390 -1218
rect 265 -1586 329 -1218
rect 984 -1586 1048 -1218
rect 1703 -1586 1767 -1218
<< mimcap >>
rect -1688 1560 -1288 1600
rect -1688 1240 -1648 1560
rect -1328 1240 -1288 1560
rect -1688 1200 -1288 1240
rect -969 1560 -569 1600
rect -969 1240 -929 1560
rect -609 1240 -569 1560
rect -969 1200 -569 1240
rect -250 1560 150 1600
rect -250 1240 -210 1560
rect 110 1240 150 1560
rect -250 1200 150 1240
rect 469 1560 869 1600
rect 469 1240 509 1560
rect 829 1240 869 1560
rect 469 1200 869 1240
rect 1188 1560 1588 1600
rect 1188 1240 1228 1560
rect 1548 1240 1588 1560
rect 1188 1200 1588 1240
rect -1688 860 -1288 900
rect -1688 540 -1648 860
rect -1328 540 -1288 860
rect -1688 500 -1288 540
rect -969 860 -569 900
rect -969 540 -929 860
rect -609 540 -569 860
rect -969 500 -569 540
rect -250 860 150 900
rect -250 540 -210 860
rect 110 540 150 860
rect -250 500 150 540
rect 469 860 869 900
rect 469 540 509 860
rect 829 540 869 860
rect 469 500 869 540
rect 1188 860 1588 900
rect 1188 540 1228 860
rect 1548 540 1588 860
rect 1188 500 1588 540
rect -1688 160 -1288 200
rect -1688 -160 -1648 160
rect -1328 -160 -1288 160
rect -1688 -200 -1288 -160
rect -969 160 -569 200
rect -969 -160 -929 160
rect -609 -160 -569 160
rect -969 -200 -569 -160
rect -250 160 150 200
rect -250 -160 -210 160
rect 110 -160 150 160
rect -250 -200 150 -160
rect 469 160 869 200
rect 469 -160 509 160
rect 829 -160 869 160
rect 469 -200 869 -160
rect 1188 160 1588 200
rect 1188 -160 1228 160
rect 1548 -160 1588 160
rect 1188 -200 1588 -160
rect -1688 -540 -1288 -500
rect -1688 -860 -1648 -540
rect -1328 -860 -1288 -540
rect -1688 -900 -1288 -860
rect -969 -540 -569 -500
rect -969 -860 -929 -540
rect -609 -860 -569 -540
rect -969 -900 -569 -860
rect -250 -540 150 -500
rect -250 -860 -210 -540
rect 110 -860 150 -540
rect -250 -900 150 -860
rect 469 -540 869 -500
rect 469 -860 509 -540
rect 829 -860 869 -540
rect 469 -900 869 -860
rect 1188 -540 1588 -500
rect 1188 -860 1228 -540
rect 1548 -860 1588 -540
rect 1188 -900 1588 -860
rect -1688 -1240 -1288 -1200
rect -1688 -1560 -1648 -1240
rect -1328 -1560 -1288 -1240
rect -1688 -1600 -1288 -1560
rect -969 -1240 -569 -1200
rect -969 -1560 -929 -1240
rect -609 -1560 -569 -1240
rect -969 -1600 -569 -1560
rect -250 -1240 150 -1200
rect -250 -1560 -210 -1240
rect 110 -1560 150 -1240
rect -250 -1600 150 -1560
rect 469 -1240 869 -1200
rect 469 -1560 509 -1240
rect 829 -1560 869 -1240
rect 469 -1600 869 -1560
rect 1188 -1240 1588 -1200
rect 1188 -1560 1228 -1240
rect 1548 -1560 1588 -1240
rect 1188 -1600 1588 -1560
<< mimcapcontact >>
rect -1648 1240 -1328 1560
rect -929 1240 -609 1560
rect -210 1240 110 1560
rect 509 1240 829 1560
rect 1228 1240 1548 1560
rect -1648 540 -1328 860
rect -929 540 -609 860
rect -210 540 110 860
rect 509 540 829 860
rect 1228 540 1548 860
rect -1648 -160 -1328 160
rect -929 -160 -609 160
rect -210 -160 110 160
rect 509 -160 829 160
rect 1228 -160 1548 160
rect -1648 -860 -1328 -540
rect -929 -860 -609 -540
rect -210 -860 110 -540
rect 509 -860 829 -540
rect 1228 -860 1548 -540
rect -1648 -1560 -1328 -1240
rect -929 -1560 -609 -1240
rect -210 -1560 110 -1240
rect 509 -1560 829 -1240
rect 1228 -1560 1548 -1240
<< metal4 >>
rect -1189 1584 -1093 1600
rect -1649 1560 -1327 1561
rect -1649 1240 -1648 1560
rect -1328 1240 -1327 1560
rect -1649 1239 -1327 1240
rect -1189 1212 -1173 1584
rect -1109 1212 -1093 1584
rect -470 1582 -374 1598
rect -930 1560 -608 1561
rect -930 1240 -929 1560
rect -609 1240 -608 1560
rect -930 1239 -608 1240
rect -1189 1196 -1093 1212
rect -470 1212 -454 1582
rect -390 1212 -374 1582
rect 249 1582 345 1598
rect -211 1560 111 1561
rect -211 1240 -210 1560
rect 110 1240 111 1560
rect -211 1239 111 1240
rect -470 1196 -374 1212
rect 249 1212 265 1582
rect 329 1212 345 1582
rect 968 1582 1064 1598
rect 508 1560 830 1561
rect 508 1240 509 1560
rect 829 1240 830 1560
rect 508 1239 830 1240
rect 249 1196 345 1212
rect 968 1212 984 1582
rect 1048 1212 1064 1582
rect 1687 1582 1783 1598
rect 1227 1560 1549 1561
rect 1227 1240 1228 1560
rect 1548 1240 1549 1560
rect 1227 1239 1549 1240
rect 968 1196 1064 1212
rect 1687 1212 1703 1582
rect 1767 1212 1783 1582
rect 1687 1196 1783 1212
rect -1189 882 -1093 898
rect -1649 860 -1327 861
rect -1649 540 -1648 860
rect -1328 540 -1327 860
rect -1649 539 -1327 540
rect -1189 514 -1173 882
rect -1109 514 -1093 882
rect -470 882 -374 898
rect -930 860 -608 861
rect -930 540 -929 860
rect -609 540 -608 860
rect -930 539 -608 540
rect -1189 494 -1093 514
rect -470 514 -454 882
rect -390 514 -374 882
rect 249 882 345 898
rect -211 860 111 861
rect -211 540 -210 860
rect 110 540 111 860
rect -211 539 111 540
rect -470 494 -374 514
rect 249 514 265 882
rect 329 514 345 882
rect 968 882 1064 898
rect 508 860 830 861
rect 508 540 509 860
rect 829 540 830 860
rect 508 539 830 540
rect 249 494 345 514
rect 968 514 984 882
rect 1048 514 1064 882
rect 1687 882 1783 898
rect 1227 860 1549 861
rect 1227 540 1228 860
rect 1548 540 1549 860
rect 1227 539 1549 540
rect 968 494 1064 514
rect 1687 514 1703 882
rect 1767 514 1783 882
rect 1687 494 1783 514
rect -1189 182 -1093 198
rect -1649 160 -1327 161
rect -1649 -160 -1648 160
rect -1328 -160 -1327 160
rect -1649 -161 -1327 -160
rect -1189 -186 -1173 182
rect -1109 -186 -1093 182
rect -470 182 -374 198
rect -930 160 -608 161
rect -930 -160 -929 160
rect -609 -160 -608 160
rect -930 -161 -608 -160
rect -1189 -204 -1093 -186
rect -470 -186 -454 182
rect -390 -186 -374 182
rect 249 182 345 198
rect -211 160 111 161
rect -211 -160 -210 160
rect 110 -160 111 160
rect -211 -161 111 -160
rect -470 -204 -374 -186
rect 249 -186 265 182
rect 329 -186 345 182
rect 968 182 1064 198
rect 508 160 830 161
rect 508 -160 509 160
rect 829 -160 830 160
rect 508 -161 830 -160
rect 249 -204 345 -186
rect 968 -186 984 182
rect 1048 -186 1064 182
rect 1687 182 1783 198
rect 1227 160 1549 161
rect 1227 -160 1228 160
rect 1548 -160 1549 160
rect 1227 -161 1549 -160
rect 968 -204 1064 -186
rect 1687 -186 1703 182
rect 1767 -186 1783 182
rect 1687 -204 1783 -186
rect -1189 -518 -1093 -502
rect -1649 -540 -1327 -539
rect -1649 -860 -1648 -540
rect -1328 -860 -1327 -540
rect -1649 -861 -1327 -860
rect -1189 -886 -1173 -518
rect -1109 -886 -1093 -518
rect -470 -518 -374 -502
rect -930 -540 -608 -539
rect -930 -860 -929 -540
rect -609 -860 -608 -540
rect -930 -861 -608 -860
rect -1189 -904 -1093 -886
rect -470 -886 -454 -518
rect -390 -886 -374 -518
rect 249 -518 345 -502
rect -211 -540 111 -539
rect -211 -860 -210 -540
rect 110 -860 111 -540
rect -211 -861 111 -860
rect -470 -904 -374 -886
rect 249 -886 265 -518
rect 329 -886 345 -518
rect 968 -518 1064 -502
rect 508 -540 830 -539
rect 508 -860 509 -540
rect 829 -860 830 -540
rect 508 -861 830 -860
rect 249 -904 345 -886
rect 968 -886 984 -518
rect 1048 -886 1064 -518
rect 1687 -518 1783 -502
rect 1227 -540 1549 -539
rect 1227 -860 1228 -540
rect 1548 -860 1549 -540
rect 1227 -861 1549 -860
rect 968 -904 1064 -886
rect 1687 -886 1703 -518
rect 1767 -886 1783 -518
rect 1687 -904 1783 -886
rect -1189 -1218 -1093 -1202
rect -1649 -1240 -1327 -1239
rect -1649 -1560 -1648 -1240
rect -1328 -1560 -1327 -1240
rect -1649 -1561 -1327 -1560
rect -1189 -1586 -1173 -1218
rect -1109 -1586 -1093 -1218
rect -470 -1218 -374 -1202
rect -930 -1240 -608 -1239
rect -930 -1560 -929 -1240
rect -609 -1560 -608 -1240
rect -930 -1561 -608 -1560
rect -1189 -1604 -1093 -1586
rect -470 -1586 -454 -1218
rect -390 -1586 -374 -1218
rect 249 -1218 345 -1202
rect -211 -1240 111 -1239
rect -211 -1560 -210 -1240
rect 110 -1560 111 -1240
rect -211 -1561 111 -1560
rect -470 -1604 -374 -1586
rect 249 -1586 265 -1218
rect 329 -1586 345 -1218
rect 968 -1218 1064 -1202
rect 508 -1240 830 -1239
rect 508 -1560 509 -1240
rect 829 -1560 830 -1240
rect 508 -1561 830 -1560
rect 249 -1604 345 -1586
rect 968 -1586 984 -1218
rect 1048 -1586 1064 -1218
rect 1687 -1218 1783 -1202
rect 1227 -1240 1549 -1239
rect 1227 -1560 1228 -1240
rect 1548 -1560 1549 -1240
rect 1227 -1561 1549 -1560
rect 968 -1604 1064 -1586
rect 1687 -1586 1703 -1218
rect 1767 -1586 1783 -1218
rect 1687 -1604 1783 -1586
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 1088 1100 1688 1700
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 5 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 0 tconnect 0 ccov 100
string library sky130
<< end >>

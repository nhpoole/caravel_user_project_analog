magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nwell >>
rect -6071 -700 6071 700
<< pmos >>
rect -5977 -600 -5177 600
rect -5119 -600 -4319 600
rect -4261 -600 -3461 600
rect -3403 -600 -2603 600
rect -2545 -600 -1745 600
rect -1687 -600 -887 600
rect -829 -600 -29 600
rect 29 -600 829 600
rect 887 -600 1687 600
rect 1745 -600 2545 600
rect 2603 -600 3403 600
rect 3461 -600 4261 600
rect 4319 -600 5119 600
rect 5177 -600 5977 600
<< pdiff >>
rect -6035 588 -5977 600
rect -6035 -588 -6023 588
rect -5989 -588 -5977 588
rect -6035 -600 -5977 -588
rect -5177 588 -5119 600
rect -5177 -588 -5165 588
rect -5131 -588 -5119 588
rect -5177 -600 -5119 -588
rect -4319 588 -4261 600
rect -4319 -588 -4307 588
rect -4273 -588 -4261 588
rect -4319 -600 -4261 -588
rect -3461 588 -3403 600
rect -3461 -588 -3449 588
rect -3415 -588 -3403 588
rect -3461 -600 -3403 -588
rect -2603 588 -2545 600
rect -2603 -588 -2591 588
rect -2557 -588 -2545 588
rect -2603 -600 -2545 -588
rect -1745 588 -1687 600
rect -1745 -588 -1733 588
rect -1699 -588 -1687 588
rect -1745 -600 -1687 -588
rect -887 588 -829 600
rect -887 -588 -875 588
rect -841 -588 -829 588
rect -887 -600 -829 -588
rect -29 588 29 600
rect -29 -588 -17 588
rect 17 -588 29 588
rect -29 -600 29 -588
rect 829 588 887 600
rect 829 -588 841 588
rect 875 -588 887 588
rect 829 -600 887 -588
rect 1687 588 1745 600
rect 1687 -588 1699 588
rect 1733 -588 1745 588
rect 1687 -600 1745 -588
rect 2545 588 2603 600
rect 2545 -588 2557 588
rect 2591 -588 2603 588
rect 2545 -600 2603 -588
rect 3403 588 3461 600
rect 3403 -588 3415 588
rect 3449 -588 3461 588
rect 3403 -600 3461 -588
rect 4261 588 4319 600
rect 4261 -588 4273 588
rect 4307 -588 4319 588
rect 4261 -600 4319 -588
rect 5119 588 5177 600
rect 5119 -588 5131 588
rect 5165 -588 5177 588
rect 5119 -600 5177 -588
rect 5977 588 6035 600
rect 5977 -588 5989 588
rect 6023 -588 6035 588
rect 5977 -600 6035 -588
<< pdiffc >>
rect -6023 -588 -5989 588
rect -5165 -588 -5131 588
rect -4307 -588 -4273 588
rect -3449 -588 -3415 588
rect -2591 -588 -2557 588
rect -1733 -588 -1699 588
rect -875 -588 -841 588
rect -17 -588 17 588
rect 841 -588 875 588
rect 1699 -588 1733 588
rect 2557 -588 2591 588
rect 3415 -588 3449 588
rect 4273 -588 4307 588
rect 5131 -588 5165 588
rect 5989 -588 6023 588
<< poly >>
rect -5823 681 -5331 697
rect -5823 664 -5807 681
rect -5977 647 -5807 664
rect -5347 664 -5331 681
rect -4965 681 -4473 697
rect -4965 664 -4949 681
rect -5347 647 -5177 664
rect -5977 600 -5177 647
rect -5119 647 -4949 664
rect -4489 664 -4473 681
rect -4107 681 -3615 697
rect -4107 664 -4091 681
rect -4489 647 -4319 664
rect -5119 600 -4319 647
rect -4261 647 -4091 664
rect -3631 664 -3615 681
rect -3249 681 -2757 697
rect -3249 664 -3233 681
rect -3631 647 -3461 664
rect -4261 600 -3461 647
rect -3403 647 -3233 664
rect -2773 664 -2757 681
rect -2391 681 -1899 697
rect -2391 664 -2375 681
rect -2773 647 -2603 664
rect -3403 600 -2603 647
rect -2545 647 -2375 664
rect -1915 664 -1899 681
rect -1533 681 -1041 697
rect -1533 664 -1517 681
rect -1915 647 -1745 664
rect -2545 600 -1745 647
rect -1687 647 -1517 664
rect -1057 664 -1041 681
rect -675 681 -183 697
rect -675 664 -659 681
rect -1057 647 -887 664
rect -1687 600 -887 647
rect -829 647 -659 664
rect -199 664 -183 681
rect 183 681 675 697
rect 183 664 199 681
rect -199 647 -29 664
rect -829 600 -29 647
rect 29 647 199 664
rect 659 664 675 681
rect 1041 681 1533 697
rect 1041 664 1057 681
rect 659 647 829 664
rect 29 600 829 647
rect 887 647 1057 664
rect 1517 664 1533 681
rect 1899 681 2391 697
rect 1899 664 1915 681
rect 1517 647 1687 664
rect 887 600 1687 647
rect 1745 647 1915 664
rect 2375 664 2391 681
rect 2757 681 3249 697
rect 2757 664 2773 681
rect 2375 647 2545 664
rect 1745 600 2545 647
rect 2603 647 2773 664
rect 3233 664 3249 681
rect 3615 681 4107 697
rect 3615 664 3631 681
rect 3233 647 3403 664
rect 2603 600 3403 647
rect 3461 647 3631 664
rect 4091 664 4107 681
rect 4473 681 4965 697
rect 4473 664 4489 681
rect 4091 647 4261 664
rect 3461 600 4261 647
rect 4319 647 4489 664
rect 4949 664 4965 681
rect 5331 681 5823 697
rect 5331 664 5347 681
rect 4949 647 5119 664
rect 4319 600 5119 647
rect 5177 647 5347 664
rect 5807 664 5823 681
rect 5807 647 5977 664
rect 5177 600 5977 647
rect -5977 -647 -5177 -600
rect -5977 -664 -5807 -647
rect -5823 -681 -5807 -664
rect -5347 -664 -5177 -647
rect -5119 -647 -4319 -600
rect -5119 -664 -4949 -647
rect -5347 -681 -5331 -664
rect -5823 -697 -5331 -681
rect -4965 -681 -4949 -664
rect -4489 -664 -4319 -647
rect -4261 -647 -3461 -600
rect -4261 -664 -4091 -647
rect -4489 -681 -4473 -664
rect -4965 -697 -4473 -681
rect -4107 -681 -4091 -664
rect -3631 -664 -3461 -647
rect -3403 -647 -2603 -600
rect -3403 -664 -3233 -647
rect -3631 -681 -3615 -664
rect -4107 -697 -3615 -681
rect -3249 -681 -3233 -664
rect -2773 -664 -2603 -647
rect -2545 -647 -1745 -600
rect -2545 -664 -2375 -647
rect -2773 -681 -2757 -664
rect -3249 -697 -2757 -681
rect -2391 -681 -2375 -664
rect -1915 -664 -1745 -647
rect -1687 -647 -887 -600
rect -1687 -664 -1517 -647
rect -1915 -681 -1899 -664
rect -2391 -697 -1899 -681
rect -1533 -681 -1517 -664
rect -1057 -664 -887 -647
rect -829 -647 -29 -600
rect -829 -664 -659 -647
rect -1057 -681 -1041 -664
rect -1533 -697 -1041 -681
rect -675 -681 -659 -664
rect -199 -664 -29 -647
rect 29 -647 829 -600
rect 29 -664 199 -647
rect -199 -681 -183 -664
rect -675 -697 -183 -681
rect 183 -681 199 -664
rect 659 -664 829 -647
rect 887 -647 1687 -600
rect 887 -664 1057 -647
rect 659 -681 675 -664
rect 183 -697 675 -681
rect 1041 -681 1057 -664
rect 1517 -664 1687 -647
rect 1745 -647 2545 -600
rect 1745 -664 1915 -647
rect 1517 -681 1533 -664
rect 1041 -697 1533 -681
rect 1899 -681 1915 -664
rect 2375 -664 2545 -647
rect 2603 -647 3403 -600
rect 2603 -664 2773 -647
rect 2375 -681 2391 -664
rect 1899 -697 2391 -681
rect 2757 -681 2773 -664
rect 3233 -664 3403 -647
rect 3461 -647 4261 -600
rect 3461 -664 3631 -647
rect 3233 -681 3249 -664
rect 2757 -697 3249 -681
rect 3615 -681 3631 -664
rect 4091 -664 4261 -647
rect 4319 -647 5119 -600
rect 4319 -664 4489 -647
rect 4091 -681 4107 -664
rect 3615 -697 4107 -681
rect 4473 -681 4489 -664
rect 4949 -664 5119 -647
rect 5177 -647 5977 -600
rect 5177 -664 5347 -647
rect 4949 -681 4965 -664
rect 4473 -697 4965 -681
rect 5331 -681 5347 -664
rect 5807 -664 5977 -647
rect 5807 -681 5823 -664
rect 5331 -697 5823 -681
<< polycont >>
rect -5807 647 -5347 681
rect -4949 647 -4489 681
rect -4091 647 -3631 681
rect -3233 647 -2773 681
rect -2375 647 -1915 681
rect -1517 647 -1057 681
rect -659 647 -199 681
rect 199 647 659 681
rect 1057 647 1517 681
rect 1915 647 2375 681
rect 2773 647 3233 681
rect 3631 647 4091 681
rect 4489 647 4949 681
rect 5347 647 5807 681
rect -5807 -681 -5347 -647
rect -4949 -681 -4489 -647
rect -4091 -681 -3631 -647
rect -3233 -681 -2773 -647
rect -2375 -681 -1915 -647
rect -1517 -681 -1057 -647
rect -659 -681 -199 -647
rect 199 -681 659 -647
rect 1057 -681 1517 -647
rect 1915 -681 2375 -647
rect 2773 -681 3233 -647
rect 3631 -681 4091 -647
rect 4489 -681 4949 -647
rect 5347 -681 5807 -647
<< locali >>
rect -5823 647 -5807 681
rect -5347 647 -5331 681
rect -4965 647 -4949 681
rect -4489 647 -4473 681
rect -4107 647 -4091 681
rect -3631 647 -3615 681
rect -3249 647 -3233 681
rect -2773 647 -2757 681
rect -2391 647 -2375 681
rect -1915 647 -1899 681
rect -1533 647 -1517 681
rect -1057 647 -1041 681
rect -675 647 -659 681
rect -199 647 -183 681
rect 183 647 199 681
rect 659 647 675 681
rect 1041 647 1057 681
rect 1517 647 1533 681
rect 1899 647 1915 681
rect 2375 647 2391 681
rect 2757 647 2773 681
rect 3233 647 3249 681
rect 3615 647 3631 681
rect 4091 647 4107 681
rect 4473 647 4489 681
rect 4949 647 4965 681
rect 5331 647 5347 681
rect 5807 647 5823 681
rect -6023 588 -5989 604
rect -6023 -604 -5989 -588
rect -5165 588 -5131 604
rect -5165 -604 -5131 -588
rect -4307 588 -4273 604
rect -4307 -604 -4273 -588
rect -3449 588 -3415 604
rect -3449 -604 -3415 -588
rect -2591 588 -2557 604
rect -2591 -604 -2557 -588
rect -1733 588 -1699 604
rect -1733 -604 -1699 -588
rect -875 588 -841 604
rect -875 -604 -841 -588
rect -17 588 17 604
rect -17 -604 17 -588
rect 841 588 875 604
rect 841 -604 875 -588
rect 1699 588 1733 604
rect 1699 -604 1733 -588
rect 2557 588 2591 604
rect 2557 -604 2591 -588
rect 3415 588 3449 604
rect 3415 -604 3449 -588
rect 4273 588 4307 604
rect 4273 -604 4307 -588
rect 5131 588 5165 604
rect 5131 -604 5165 -588
rect 5989 588 6023 604
rect 5989 -604 6023 -588
rect -5823 -681 -5807 -647
rect -5347 -681 -5331 -647
rect -4965 -681 -4949 -647
rect -4489 -681 -4473 -647
rect -4107 -681 -4091 -647
rect -3631 -681 -3615 -647
rect -3249 -681 -3233 -647
rect -2773 -681 -2757 -647
rect -2391 -681 -2375 -647
rect -1915 -681 -1899 -647
rect -1533 -681 -1517 -647
rect -1057 -681 -1041 -647
rect -675 -681 -659 -647
rect -199 -681 -183 -647
rect 183 -681 199 -647
rect 659 -681 675 -647
rect 1041 -681 1057 -647
rect 1517 -681 1533 -647
rect 1899 -681 1915 -647
rect 2375 -681 2391 -647
rect 2757 -681 2773 -647
rect 3233 -681 3249 -647
rect 3615 -681 3631 -647
rect 4091 -681 4107 -647
rect 4473 -681 4489 -647
rect 4949 -681 4965 -647
rect 5331 -681 5347 -647
rect 5807 -681 5823 -647
<< viali >>
rect -5769 647 -5385 681
rect -4911 647 -4527 681
rect -4053 647 -3669 681
rect -3195 647 -2811 681
rect -2337 647 -1953 681
rect -1479 647 -1095 681
rect -621 647 -237 681
rect 237 647 621 681
rect 1095 647 1479 681
rect 1953 647 2337 681
rect 2811 647 3195 681
rect 3669 647 4053 681
rect 4527 647 4911 681
rect 5385 647 5769 681
rect -6023 -588 -5989 588
rect -5165 -588 -5131 588
rect -4307 -588 -4273 588
rect -3449 -588 -3415 588
rect -2591 -588 -2557 588
rect -1733 -588 -1699 588
rect -875 -588 -841 588
rect -17 -588 17 588
rect 841 -588 875 588
rect 1699 -588 1733 588
rect 2557 -588 2591 588
rect 3415 -588 3449 588
rect 4273 -588 4307 588
rect 5131 -588 5165 588
rect 5989 -588 6023 588
rect -5769 -681 -5385 -647
rect -4911 -681 -4527 -647
rect -4053 -681 -3669 -647
rect -3195 -681 -2811 -647
rect -2337 -681 -1953 -647
rect -1479 -681 -1095 -647
rect -621 -681 -237 -647
rect 237 -681 621 -647
rect 1095 -681 1479 -647
rect 1953 -681 2337 -647
rect 2811 -681 3195 -647
rect 3669 -681 4053 -647
rect 4527 -681 4911 -647
rect 5385 -681 5769 -647
<< metal1 >>
rect -5781 681 -5373 687
rect -5781 647 -5769 681
rect -5385 647 -5373 681
rect -5781 641 -5373 647
rect -4923 681 -4515 687
rect -4923 647 -4911 681
rect -4527 647 -4515 681
rect -4923 641 -4515 647
rect -4065 681 -3657 687
rect -4065 647 -4053 681
rect -3669 647 -3657 681
rect -4065 641 -3657 647
rect -3207 681 -2799 687
rect -3207 647 -3195 681
rect -2811 647 -2799 681
rect -3207 641 -2799 647
rect -2349 681 -1941 687
rect -2349 647 -2337 681
rect -1953 647 -1941 681
rect -2349 641 -1941 647
rect -1491 681 -1083 687
rect -1491 647 -1479 681
rect -1095 647 -1083 681
rect -1491 641 -1083 647
rect -633 681 -225 687
rect -633 647 -621 681
rect -237 647 -225 681
rect -633 641 -225 647
rect 225 681 633 687
rect 225 647 237 681
rect 621 647 633 681
rect 225 641 633 647
rect 1083 681 1491 687
rect 1083 647 1095 681
rect 1479 647 1491 681
rect 1083 641 1491 647
rect 1941 681 2349 687
rect 1941 647 1953 681
rect 2337 647 2349 681
rect 1941 641 2349 647
rect 2799 681 3207 687
rect 2799 647 2811 681
rect 3195 647 3207 681
rect 2799 641 3207 647
rect 3657 681 4065 687
rect 3657 647 3669 681
rect 4053 647 4065 681
rect 3657 641 4065 647
rect 4515 681 4923 687
rect 4515 647 4527 681
rect 4911 647 4923 681
rect 4515 641 4923 647
rect 5373 681 5781 687
rect 5373 647 5385 681
rect 5769 647 5781 681
rect 5373 641 5781 647
rect -6029 588 -5983 600
rect -6029 -588 -6023 588
rect -5989 -588 -5983 588
rect -6029 -600 -5983 -588
rect -5171 588 -5125 600
rect -5171 -588 -5165 588
rect -5131 -588 -5125 588
rect -5171 -600 -5125 -588
rect -4313 588 -4267 600
rect -4313 -588 -4307 588
rect -4273 -588 -4267 588
rect -4313 -600 -4267 -588
rect -3455 588 -3409 600
rect -3455 -588 -3449 588
rect -3415 -588 -3409 588
rect -3455 -600 -3409 -588
rect -2597 588 -2551 600
rect -2597 -588 -2591 588
rect -2557 -588 -2551 588
rect -2597 -600 -2551 -588
rect -1739 588 -1693 600
rect -1739 -588 -1733 588
rect -1699 -588 -1693 588
rect -1739 -600 -1693 -588
rect -881 588 -835 600
rect -881 -588 -875 588
rect -841 -588 -835 588
rect -881 -600 -835 -588
rect -23 588 23 600
rect -23 -588 -17 588
rect 17 -588 23 588
rect -23 -600 23 -588
rect 835 588 881 600
rect 835 -588 841 588
rect 875 -588 881 588
rect 835 -600 881 -588
rect 1693 588 1739 600
rect 1693 -588 1699 588
rect 1733 -588 1739 588
rect 1693 -600 1739 -588
rect 2551 588 2597 600
rect 2551 -588 2557 588
rect 2591 -588 2597 588
rect 2551 -600 2597 -588
rect 3409 588 3455 600
rect 3409 -588 3415 588
rect 3449 -588 3455 588
rect 3409 -600 3455 -588
rect 4267 588 4313 600
rect 4267 -588 4273 588
rect 4307 -588 4313 588
rect 4267 -600 4313 -588
rect 5125 588 5171 600
rect 5125 -588 5131 588
rect 5165 -588 5171 588
rect 5125 -600 5171 -588
rect 5983 588 6029 600
rect 5983 -588 5989 588
rect 6023 -588 6029 588
rect 5983 -600 6029 -588
rect -5781 -647 -5373 -641
rect -5781 -681 -5769 -647
rect -5385 -681 -5373 -647
rect -5781 -687 -5373 -681
rect -4923 -647 -4515 -641
rect -4923 -681 -4911 -647
rect -4527 -681 -4515 -647
rect -4923 -687 -4515 -681
rect -4065 -647 -3657 -641
rect -4065 -681 -4053 -647
rect -3669 -681 -3657 -647
rect -4065 -687 -3657 -681
rect -3207 -647 -2799 -641
rect -3207 -681 -3195 -647
rect -2811 -681 -2799 -647
rect -3207 -687 -2799 -681
rect -2349 -647 -1941 -641
rect -2349 -681 -2337 -647
rect -1953 -681 -1941 -647
rect -2349 -687 -1941 -681
rect -1491 -647 -1083 -641
rect -1491 -681 -1479 -647
rect -1095 -681 -1083 -647
rect -1491 -687 -1083 -681
rect -633 -647 -225 -641
rect -633 -681 -621 -647
rect -237 -681 -225 -647
rect -633 -687 -225 -681
rect 225 -647 633 -641
rect 225 -681 237 -647
rect 621 -681 633 -647
rect 225 -687 633 -681
rect 1083 -647 1491 -641
rect 1083 -681 1095 -647
rect 1479 -681 1491 -647
rect 1083 -687 1491 -681
rect 1941 -647 2349 -641
rect 1941 -681 1953 -647
rect 2337 -681 2349 -647
rect 1941 -687 2349 -681
rect 2799 -647 3207 -641
rect 2799 -681 2811 -647
rect 3195 -681 3207 -647
rect 2799 -687 3207 -681
rect 3657 -647 4065 -641
rect 3657 -681 3669 -647
rect 4053 -681 4065 -647
rect 3657 -687 4065 -681
rect 4515 -647 4923 -641
rect 4515 -681 4527 -647
rect 4911 -681 4923 -647
rect 4515 -687 4923 -681
rect 5373 -647 5781 -641
rect 5373 -681 5385 -647
rect 5769 -681 5781 -647
rect 5373 -687 5781 -681
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 6 l 4 m 1 nf 14 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nwell >>
rect -5058 4282 5458 10358
<< pwell >>
rect -5058 1752 5458 4118
<< psubdiff >>
rect -5022 4142 -4860 4242
rect 5260 4142 5422 4242
rect -5022 4080 -4922 4142
rect -5022 1878 -4922 1940
rect 5322 4080 5422 4142
rect 5322 1878 5422 1940
rect -5022 1778 -4860 1878
rect 5260 1778 5422 1878
<< nsubdiff >>
rect -5022 10222 -4860 10322
rect 5260 10222 5422 10322
rect -5022 10160 -4922 10222
rect -5022 4578 -4922 4640
rect 5322 10160 5422 10222
rect 5322 4578 5422 4640
rect -5022 4478 -4860 4578
rect 5260 4478 5422 4578
<< psubdiffcont >>
rect -4860 4142 5260 4242
rect -5022 1940 -4922 4080
rect 5322 1940 5422 4080
rect -4860 1778 5260 1878
<< nsubdiffcont >>
rect -4860 10222 5260 10322
rect -5022 4640 -4922 10160
rect 5322 4640 5422 10160
rect -4860 4478 5260 4578
<< locali >>
rect -5022 10160 -4922 10322
rect 5322 10160 5422 10322
rect -158 7106 302 7112
rect -158 7058 -152 7106
rect -104 7058 302 7106
rect -158 7052 302 7058
rect -5022 4478 -4922 4640
rect 5322 4478 5422 4640
rect -5022 4080 -4922 4242
rect -5022 1778 -4922 1940
rect 5322 4080 5422 4242
rect 5322 1778 5422 1940
<< viali >>
rect -4922 10222 -4860 10322
rect -4860 10222 5260 10322
rect 5260 10222 5322 10322
rect -5022 4760 -4922 9932
rect -152 7058 -104 7106
rect 302 7052 362 7112
rect 5322 4760 5422 9932
rect -4922 4478 -4860 4578
rect -4860 4478 5260 4578
rect 5260 4478 5322 4578
rect -4922 4142 -4860 4242
rect -4860 4142 5260 4242
rect 5260 4142 5322 4242
rect -5022 2008 -4922 4012
rect 5322 2008 5422 4012
rect -4922 1778 -4860 1878
rect -4860 1778 5260 1878
rect 5260 1778 5322 1878
<< metal1 >>
rect -5028 10322 5428 10328
rect -5028 10222 -4922 10322
rect 5322 10222 5428 10322
rect -5028 10216 5428 10222
rect -5028 9932 -4916 10216
rect -5028 4760 -5022 9932
rect -4922 7110 -4916 9932
rect -4316 9916 -4306 10216
rect 4706 9916 4716 10216
rect 5316 9932 5428 10216
rect -4078 9742 4278 9756
rect -4078 9656 -4064 9742
rect -3968 9656 -3464 9742
rect -3368 9656 -2864 9742
rect -2768 9656 -2264 9742
rect -2168 9656 -1664 9742
rect -1568 9656 -1064 9742
rect -968 9656 -464 9742
rect -368 9656 136 9742
rect 232 9656 736 9742
rect 832 9656 1336 9742
rect 1432 9656 1936 9742
rect 2032 9656 2536 9742
rect 2632 9656 3136 9742
rect 3232 9656 3736 9742
rect 3832 9656 4156 9742
rect 4252 9656 4278 9742
rect -4078 9646 4278 9656
rect -4050 8826 -3990 9646
rect -3818 8918 -3758 9646
rect -3592 8794 -3532 9646
rect -2676 9392 2882 9452
rect -3366 9024 -3360 9084
rect -3300 9024 -3294 9084
rect -2910 9024 -2904 9084
rect -2844 9024 -2838 9084
rect -3360 8916 -3300 9024
rect -2904 8918 -2844 9024
rect -2676 8800 -2616 9392
rect -1760 9258 1962 9318
rect -2450 9024 -2444 9084
rect -2384 9024 -2378 9084
rect -1994 9024 -1988 9084
rect -1928 9024 -1922 9084
rect -2444 8912 -2384 9024
rect -1988 8918 -1928 9024
rect -1760 8798 -1700 9258
rect -844 9134 1046 9194
rect -1536 9024 -1530 9084
rect -1470 9024 -1464 9084
rect -1072 9024 -1066 9084
rect -1006 9024 -1000 9084
rect -1530 8918 -1470 9024
rect -1066 8914 -1006 9024
rect -844 8780 -784 9134
rect -622 9024 -616 9084
rect -556 9024 -550 9084
rect -166 9024 -160 9084
rect -100 9024 -94 9084
rect 302 9024 308 9084
rect 368 9024 374 9084
rect 760 9024 766 9084
rect 826 9024 832 9084
rect -616 8920 -556 9024
rect -160 8920 -100 9024
rect 308 8920 368 9024
rect 766 8924 826 9024
rect 986 8814 1046 9134
rect 1216 9024 1222 9084
rect 1282 9024 1288 9084
rect 1672 9024 1678 9084
rect 1738 9024 1744 9084
rect 1222 8918 1282 9024
rect 1678 8918 1738 9024
rect 1902 8800 1962 9258
rect 2128 9024 2134 9084
rect 2194 9024 2200 9084
rect 2584 9024 2590 9084
rect 2650 9024 2656 9084
rect 2134 8918 2194 9024
rect 2590 8922 2650 9024
rect 2822 8802 2882 9392
rect 3042 9024 3048 9084
rect 3108 9024 3114 9084
rect 3502 9024 3508 9084
rect 3568 9024 3574 9084
rect 3048 8918 3108 9024
rect 3508 8914 3568 9024
rect 3738 8782 3798 9646
rect 3968 8916 4028 9646
rect 4196 8788 4256 9646
rect -4048 7110 -3988 7342
rect -3820 7110 -3760 7226
rect -3594 7110 -3534 7326
rect -3364 7110 -3304 7218
rect -4922 7050 -3534 7110
rect -3370 7050 -3364 7110
rect -3304 7050 -3298 7110
rect -4922 6678 -4916 7050
rect -4048 6678 -3988 7050
rect -4922 6618 -3988 6678
rect -3136 6630 -3076 7366
rect -2908 7110 -2848 7216
rect -2448 7110 -2388 7222
rect -2914 7050 -2908 7110
rect -2848 7050 -2842 7110
rect -2454 7050 -2448 7110
rect -2388 7050 -2382 7110
rect -2218 6760 -2158 7360
rect -1992 7110 -1932 7216
rect -1534 7110 -1474 7216
rect -1998 7050 -1992 7110
rect -1932 7050 -1926 7110
rect -1540 7050 -1534 7110
rect -1474 7050 -1468 7110
rect -1310 6886 -1250 7354
rect -1070 7110 -1010 7220
rect -616 7110 -556 7222
rect -1076 7050 -1070 7110
rect -1010 7050 -1004 7110
rect -622 7050 -616 7110
rect -556 7050 -550 7110
rect -386 7002 -326 7362
rect -158 7112 -98 7220
rect 76 7122 136 7304
rect -164 7110 -92 7112
rect -164 7050 -158 7110
rect -98 7050 -92 7110
rect 302 7118 362 7228
rect 76 7056 136 7062
rect 290 7112 374 7118
rect 290 7050 302 7112
rect 362 7050 374 7112
rect 290 7046 374 7050
rect 532 7002 592 7310
rect 758 7110 818 7222
rect 1218 7110 1278 7216
rect 752 7050 758 7110
rect 818 7050 824 7110
rect 1212 7050 1218 7110
rect 1278 7050 1284 7110
rect -386 6942 592 7002
rect 1446 6886 1506 7314
rect 1674 7110 1734 7216
rect 2130 7110 2190 7216
rect 1668 7050 1674 7110
rect 1734 7050 1740 7110
rect 2124 7050 2130 7110
rect 2190 7050 2196 7110
rect -1310 6826 1506 6886
rect 2366 6760 2426 7350
rect 2586 7110 2646 7212
rect 3044 7110 3104 7216
rect 2580 7050 2586 7110
rect 2646 7050 2652 7110
rect 3038 7050 3044 7110
rect 3104 7050 3110 7110
rect -2218 6700 2426 6760
rect 3280 6630 3340 7342
rect 3504 7110 3564 7220
rect 3498 7050 3504 7110
rect 3564 7050 3570 7110
rect 3734 7108 3794 7344
rect 3966 7108 4026 7224
rect 4192 7108 4252 7326
rect 5316 7108 5322 9932
rect 3734 7048 5322 7108
rect -4922 4760 -4916 6618
rect -4608 6146 -4548 6618
rect -4380 6254 -4320 6618
rect -3136 6570 3340 6630
rect 4192 6614 4252 7048
rect 5316 6614 5322 7048
rect 4192 6554 5322 6614
rect -4156 6464 -4150 6524
rect -4090 6464 -4084 6524
rect -4150 6126 -4090 6464
rect -3918 6362 -654 6422
rect -3918 6250 -3858 6362
rect -3456 6266 -3396 6362
rect -3002 6260 -2942 6362
rect -2540 6260 -2480 6362
rect -2086 6260 -2026 6362
rect -1636 6266 -1576 6362
rect -1170 6272 -1110 6362
rect -714 6266 -654 6362
rect -258 6344 910 6404
rect -258 6254 -198 6344
rect -28 6178 32 6344
rect 392 6172 452 6344
rect 624 6254 684 6344
rect 850 6150 910 6344
rect 1076 6362 4340 6422
rect 1076 6250 1136 6362
rect 1538 6266 1598 6362
rect 1992 6260 2052 6362
rect 2454 6260 2514 6362
rect 2908 6260 2968 6362
rect 3358 6266 3418 6362
rect 3824 6272 3884 6362
rect 4280 6266 4340 6362
rect 4742 6256 4802 6554
rect 4968 6140 5028 6554
rect -5028 4584 -4916 4760
rect -4608 4584 -4548 5038
rect -4380 4584 -4320 4958
rect -3926 4850 -3866 4962
rect -3464 4850 -3404 4946
rect -3010 4850 -2950 4952
rect -2548 4850 -2488 4952
rect -2094 4850 -2034 4952
rect -1644 4850 -1584 4946
rect -1178 4850 -1118 4940
rect -722 4850 -662 4946
rect -3926 4846 -3010 4850
rect -3866 4790 -3464 4846
rect -3926 4780 -3866 4786
rect -3404 4790 -3010 4846
rect -2950 4790 -2548 4850
rect -2488 4844 -1644 4850
rect -2488 4790 -2094 4844
rect -3464 4780 -3404 4786
rect -3010 4784 -2950 4790
rect -2548 4784 -2488 4790
rect -2034 4790 -1644 4844
rect -1584 4790 -1178 4850
rect -1118 4846 -662 4850
rect -1118 4790 -722 4846
rect -1644 4784 -1584 4790
rect -1178 4784 -1118 4790
rect -2094 4778 -2034 4784
rect -722 4780 -662 4786
rect -488 4724 -428 5084
rect -494 4664 -488 4724
rect -428 4664 -422 4724
rect -258 4584 -198 4960
rect -30 4584 30 5052
rect 390 4584 450 5052
rect 618 4584 678 4956
rect 848 4584 908 5058
rect 1076 4850 1136 4962
rect 1538 4854 1598 4946
rect 1076 4846 1538 4850
rect 1136 4794 1538 4846
rect 1992 4850 2052 4952
rect 2454 4850 2514 4952
rect 2908 4850 2968 4952
rect 3358 4854 3418 4946
rect 1598 4848 3358 4850
rect 1598 4794 1992 4848
rect 1136 4790 1992 4794
rect 1538 4788 1598 4790
rect 2052 4790 2454 4848
rect 1076 4780 1136 4786
rect 1992 4782 2052 4788
rect 2514 4790 2908 4848
rect 2454 4782 2514 4788
rect 2968 4794 3358 4848
rect 3824 4850 3884 4940
rect 4280 4850 4340 4946
rect 3418 4848 4340 4850
rect 3418 4794 3824 4848
rect 2968 4790 3824 4794
rect 3358 4788 3418 4790
rect 3884 4790 4280 4848
rect 2908 4782 2968 4788
rect 3824 4782 3884 4788
rect 4280 4782 4340 4788
rect 4512 4718 4572 5024
rect 4512 4652 4572 4658
rect 4742 4584 4802 4956
rect 4970 4584 5030 5050
rect 5316 4760 5322 6554
rect 5422 4760 5428 9932
rect 5316 4584 5428 4760
rect -5028 4578 5428 4584
rect -5028 4478 -4922 4578
rect 5322 4478 5428 4578
rect -5028 4472 5428 4478
rect -5028 4242 5428 4248
rect -5028 4142 -4922 4242
rect 5322 4142 5428 4242
rect -5028 4136 5428 4142
rect -5028 4012 -4916 4136
rect -5028 2008 -5022 4012
rect -4922 2008 -4916 4012
rect -4608 3660 -4548 4136
rect -4378 3748 -4318 4136
rect -488 4044 -428 4050
rect -3920 3910 -3464 3916
rect -3932 3850 -3926 3910
rect -3866 3856 -3464 3910
rect -3404 3910 -2548 3916
rect -3404 3856 -3010 3910
rect -3866 3850 -3860 3856
rect -3926 3754 -3860 3850
rect -3920 3750 -3860 3754
rect -3464 3760 -3398 3856
rect -3016 3850 -3010 3856
rect -2950 3856 -2548 3910
rect -2488 3856 -2094 3916
rect -2034 3856 -1644 3916
rect -1584 3910 -722 3916
rect -1584 3856 -1178 3910
rect -2950 3850 -2944 3856
rect -3464 3752 -3404 3760
rect -3010 3758 -2944 3850
rect -3004 3754 -2944 3758
rect -2548 3754 -2482 3856
rect -2094 3758 -2028 3856
rect -2088 3754 -2028 3758
rect -1644 3760 -1578 3856
rect -1184 3850 -1178 3856
rect -1118 3856 -722 3910
rect -662 3856 -656 3916
rect -1118 3850 -1112 3856
rect -1178 3766 -1112 3850
rect -1644 3748 -1584 3760
rect -1178 3748 -1118 3766
rect -722 3760 -656 3856
rect -722 3758 -662 3760
rect -488 3670 -428 3984
rect -260 3752 -200 4136
rect -28 3672 32 4136
rect 392 3664 452 4136
rect 626 3752 686 4136
rect 848 3636 908 4136
rect 4506 3996 4512 4056
rect 4572 3996 4578 4056
rect 3352 3916 3358 3920
rect 1070 3856 1076 3916
rect 1136 3914 3358 3916
rect 1136 3856 1538 3914
rect 1076 3750 1140 3856
rect 1532 3854 1538 3856
rect 1598 3856 1992 3914
rect 1598 3854 1604 3856
rect 1986 3854 1992 3856
rect 2052 3856 2454 3914
rect 2052 3854 2058 3856
rect 2448 3854 2454 3856
rect 2514 3856 2908 3914
rect 2514 3854 2520 3856
rect 2902 3854 2908 3856
rect 2968 3860 3358 3914
rect 3418 3916 3424 3920
rect 3418 3860 3824 3916
rect 2968 3856 3824 3860
rect 3884 3856 4280 3916
rect 4340 3856 4346 3916
rect 2968 3854 2974 3856
rect 1538 3760 1602 3854
rect 1538 3752 1598 3760
rect 1992 3754 2056 3854
rect 2454 3754 2518 3854
rect 2908 3754 2972 3854
rect 3358 3760 3422 3856
rect 3824 3766 3888 3856
rect 1076 3746 1136 3750
rect 1992 3746 2052 3754
rect 2454 3748 2514 3754
rect 2908 3748 2968 3754
rect 3358 3752 3418 3760
rect 3824 3752 3884 3766
rect 4280 3760 4344 3856
rect 4280 3748 4340 3760
rect 4512 3658 4572 3996
rect 4752 3754 4812 4136
rect 4970 3660 5030 4136
rect 5316 4012 5428 4136
rect -4608 3308 -4548 3564
rect -4380 3308 -4320 3472
rect -4608 3248 -4320 3308
rect -4608 3012 -4548 3248
rect -4380 3082 -4320 3248
rect -4152 3004 -4092 3566
rect -3926 3368 -3866 3474
rect -3464 3368 -3404 3464
rect -3010 3368 -2950 3470
rect -2548 3368 -2488 3470
rect -2094 3368 -2034 3470
rect -1644 3368 -1584 3464
rect -1178 3368 -1118 3458
rect -722 3368 -662 3464
rect -3926 3308 -662 3368
rect -3920 3188 -656 3248
rect -3920 3082 -3860 3188
rect -3458 3092 -3398 3188
rect -3004 3086 -2944 3188
rect -2542 3086 -2482 3188
rect -2088 3086 -2028 3188
rect -1638 3092 -1578 3188
rect -1172 3098 -1112 3188
rect -716 3092 -656 3188
rect -260 3084 -200 3476
rect -4616 2476 -4556 2886
rect -4376 2476 -4316 2806
rect -3926 2700 -3866 2806
rect -3464 2700 -3404 2796
rect -3010 2700 -2950 2802
rect -2548 2700 -2488 2802
rect -2094 2700 -2034 2802
rect -1644 2700 -1584 2796
rect -1178 2700 -1118 2790
rect -722 2700 -662 2796
rect -3926 2640 -662 2700
rect -488 2476 -428 2884
rect -262 2476 -202 2808
rect -28 2476 32 3580
rect 388 3370 448 3560
rect 616 3370 676 3478
rect 848 3370 908 3568
rect 388 3310 908 3370
rect 388 2476 448 3310
rect 616 2476 676 3310
rect 848 2476 908 3310
rect 1074 3368 1134 3474
rect 1536 3368 1596 3464
rect 1990 3368 2050 3470
rect 2452 3368 2512 3470
rect 2906 3368 2966 3470
rect 3356 3368 3416 3464
rect 3822 3368 3882 3458
rect 4278 3368 4338 3464
rect 1074 3308 4338 3368
rect 4742 2476 4802 3474
rect 4968 2476 5028 3570
rect -4680 2448 5090 2476
rect -4680 2362 -4630 2448
rect -4534 2362 -4050 2448
rect -3954 2362 -3450 2448
rect -3354 2362 -2850 2448
rect -2754 2362 -2250 2448
rect -2154 2362 -1650 2448
rect -1554 2362 -1050 2448
rect -954 2362 -450 2448
rect -354 2362 150 2448
rect 246 2362 750 2448
rect 846 2362 1350 2448
rect 1446 2362 1950 2448
rect 2046 2362 2550 2448
rect 2646 2362 3150 2448
rect 3246 2362 3750 2448
rect 3846 2362 4350 2448
rect 4446 2362 4950 2448
rect 5046 2362 5090 2448
rect -4680 2332 5090 2362
rect -5028 1884 -4916 2008
rect -4316 1884 -4306 2184
rect 4706 1884 4716 2184
rect 5316 2008 5322 4012
rect 5422 2008 5428 4012
rect 5316 1884 5428 2008
rect -5028 1878 5428 1884
rect -5028 1778 -4922 1878
rect 5322 1778 5428 1878
rect -5028 1772 5428 1778
<< via1 >>
rect -4916 9916 -4316 10216
rect 4716 9916 5316 10216
rect -4064 9656 -3968 9742
rect -3464 9656 -3368 9742
rect -2864 9656 -2768 9742
rect -2264 9656 -2168 9742
rect -1664 9656 -1568 9742
rect -1064 9656 -968 9742
rect -464 9656 -368 9742
rect 136 9656 232 9742
rect 736 9656 832 9742
rect 1336 9656 1432 9742
rect 1936 9656 2032 9742
rect 2536 9656 2632 9742
rect 3136 9656 3232 9742
rect 3736 9656 3832 9742
rect 4156 9656 4252 9742
rect -3360 9024 -3300 9084
rect -2904 9024 -2844 9084
rect -2444 9024 -2384 9084
rect -1988 9024 -1928 9084
rect -1530 9024 -1470 9084
rect -1066 9024 -1006 9084
rect -616 9024 -556 9084
rect -160 9024 -100 9084
rect 308 9024 368 9084
rect 766 9024 826 9084
rect 1222 9024 1282 9084
rect 1678 9024 1738 9084
rect 2134 9024 2194 9084
rect 2590 9024 2650 9084
rect 3048 9024 3108 9084
rect 3508 9024 3568 9084
rect -3364 7050 -3304 7110
rect -2908 7050 -2848 7110
rect -2448 7050 -2388 7110
rect -1992 7050 -1932 7110
rect -1534 7050 -1474 7110
rect -1070 7050 -1010 7110
rect -616 7050 -556 7110
rect -158 7106 -98 7110
rect -158 7058 -152 7106
rect -152 7058 -104 7106
rect -104 7058 -98 7106
rect -158 7050 -98 7058
rect 76 7062 136 7122
rect 302 7052 362 7110
rect 302 7050 362 7052
rect 758 7050 818 7110
rect 1218 7050 1278 7110
rect 1674 7050 1734 7110
rect 2130 7050 2190 7110
rect 2586 7050 2646 7110
rect 3044 7050 3104 7110
rect 3504 7050 3564 7110
rect -4150 6464 -4090 6524
rect -3926 4786 -3866 4846
rect -3464 4786 -3404 4846
rect -3010 4790 -2950 4850
rect -2548 4790 -2488 4850
rect -2094 4784 -2034 4844
rect -1644 4790 -1584 4850
rect -1178 4790 -1118 4850
rect -722 4786 -662 4846
rect -488 4664 -428 4724
rect 1076 4786 1136 4846
rect 1538 4794 1598 4854
rect 1992 4788 2052 4848
rect 2454 4788 2514 4848
rect 2908 4788 2968 4848
rect 3358 4794 3418 4854
rect 3824 4788 3884 4848
rect 4280 4788 4340 4848
rect 4512 4658 4572 4718
rect -488 3984 -428 4044
rect -3926 3850 -3866 3910
rect -3464 3856 -3404 3916
rect -3010 3850 -2950 3910
rect -2548 3856 -2488 3916
rect -2094 3856 -2034 3916
rect -1644 3856 -1584 3916
rect -1178 3850 -1118 3910
rect -722 3856 -662 3916
rect 4512 3996 4572 4056
rect 1076 3856 1136 3916
rect 1538 3854 1598 3914
rect 1992 3854 2052 3914
rect 2454 3854 2514 3914
rect 2908 3854 2968 3914
rect 3358 3860 3418 3920
rect 3824 3856 3884 3916
rect 4280 3856 4340 3916
rect -4630 2362 -4534 2448
rect -4050 2362 -3954 2448
rect -3450 2362 -3354 2448
rect -2850 2362 -2754 2448
rect -2250 2362 -2154 2448
rect -1650 2362 -1554 2448
rect -1050 2362 -954 2448
rect -450 2362 -354 2448
rect 150 2362 246 2448
rect 750 2362 846 2448
rect 1350 2362 1446 2448
rect 1950 2362 2046 2448
rect 2550 2362 2646 2448
rect 3150 2362 3246 2448
rect 3750 2362 3846 2448
rect 4350 2362 4446 2448
rect 4950 2362 5046 2448
rect -4916 1884 -4316 2184
rect 4716 1884 5316 2184
<< metal2 >>
rect -4916 10216 -4316 10226
rect -4916 9906 -4316 9916
rect 4716 10216 5316 10226
rect 4716 9906 5316 9916
rect -4078 9742 4278 9756
rect -4078 9656 -4064 9742
rect -3968 9656 -3464 9742
rect -3368 9656 -2864 9742
rect -2768 9656 -2264 9742
rect -2168 9656 -1664 9742
rect -1568 9656 -1064 9742
rect -968 9656 -464 9742
rect -368 9656 136 9742
rect 232 9656 736 9742
rect 832 9656 1336 9742
rect 1432 9656 1936 9742
rect 2032 9656 2536 9742
rect 2632 9656 3136 9742
rect 3232 9656 3736 9742
rect 3832 9656 4156 9742
rect 4252 9656 4278 9742
rect -4078 9646 4278 9656
rect -3360 9084 -3300 9090
rect -2904 9084 -2844 9090
rect -2444 9084 -2384 9090
rect -1988 9084 -1928 9090
rect -1530 9084 -1470 9090
rect -1066 9084 -1006 9090
rect -616 9084 -556 9090
rect -160 9084 -100 9090
rect 308 9084 368 9090
rect 766 9084 826 9090
rect 1222 9084 1282 9090
rect 1678 9084 1738 9090
rect 2134 9084 2194 9090
rect 2590 9084 2650 9090
rect 3048 9084 3108 9090
rect 3508 9084 3568 9090
rect -3300 9024 -2904 9084
rect -2844 9024 -2444 9084
rect -2384 9024 -1988 9084
rect -1928 9024 -1530 9084
rect -1470 9024 -1066 9084
rect -1006 9024 -616 9084
rect -556 9024 -160 9084
rect -100 9024 308 9084
rect 368 9024 766 9084
rect 826 9024 1222 9084
rect 1282 9024 1678 9084
rect 1738 9024 2134 9084
rect 2194 9024 2590 9084
rect 2650 9024 3048 9084
rect 3108 9024 3508 9084
rect -3360 9018 -3300 9024
rect -2904 9018 -2844 9024
rect -2444 9018 -2384 9024
rect -1988 9018 -1928 9024
rect -1530 9018 -1470 9024
rect -1066 9018 -1006 9024
rect -616 9018 -556 9024
rect -160 9018 -100 9024
rect 308 9018 368 9024
rect 766 9018 826 9024
rect 1222 9018 1282 9024
rect 1678 9018 1738 9024
rect 2134 9018 2194 9024
rect 2590 9018 2650 9024
rect 3048 9018 3108 9024
rect 3508 9018 3568 9024
rect -3364 7110 -3304 7116
rect -2908 7110 -2848 7116
rect -2448 7110 -2388 7116
rect -1992 7110 -1932 7116
rect -1534 7110 -1474 7116
rect -1070 7110 -1010 7116
rect -616 7110 -556 7116
rect -158 7110 -98 7116
rect -3304 7050 -2908 7110
rect -2848 7050 -2448 7110
rect -2388 7050 -1992 7110
rect -1932 7050 -1534 7110
rect -1474 7050 -1070 7110
rect -1010 7050 -616 7110
rect -556 7050 -158 7110
rect 70 7062 76 7122
rect 136 7062 142 7122
rect 302 7110 362 7116
rect 758 7110 818 7116
rect 1218 7110 1278 7116
rect 1674 7110 1734 7116
rect 2130 7110 2190 7116
rect 2586 7110 2646 7116
rect 3044 7110 3104 7116
rect 3504 7110 3564 7116
rect -3364 7044 -3304 7050
rect -2908 7044 -2848 7050
rect -2448 7044 -2388 7050
rect -1992 7044 -1932 7050
rect -1534 7044 -1474 7050
rect -1070 7044 -1010 7050
rect -616 7044 -556 7050
rect -158 7044 -98 7050
rect -4150 6524 -4090 6530
rect 76 6524 136 7062
rect 362 7050 758 7110
rect 818 7050 1218 7110
rect 1278 7050 1674 7110
rect 1734 7050 2130 7110
rect 2190 7050 2586 7110
rect 2646 7050 3044 7110
rect 3104 7050 3504 7110
rect 302 7044 362 7050
rect 758 7044 818 7050
rect 1218 7044 1278 7050
rect 1674 7044 1734 7050
rect 2130 7044 2190 7050
rect 2586 7044 2646 7050
rect 3044 7044 3104 7050
rect 3504 7044 3564 7050
rect -4090 6464 136 6524
rect -4150 6458 -4090 6464
rect -3932 4786 -3926 4846
rect -3866 4786 -3860 4846
rect -3470 4786 -3464 4846
rect -3404 4786 -3398 4846
rect -3016 4790 -3010 4850
rect -2950 4790 -2944 4850
rect -2554 4790 -2548 4850
rect -2488 4790 -2482 4850
rect -3926 4392 -3866 4786
rect -3464 4392 -3404 4786
rect -3010 4392 -2950 4790
rect -2548 4392 -2488 4790
rect -2100 4784 -2094 4844
rect -2034 4784 -2028 4844
rect -1650 4790 -1644 4850
rect -1584 4790 -1578 4850
rect -1184 4790 -1178 4850
rect -1118 4790 -1112 4850
rect -2094 4392 -2034 4784
rect -1644 4392 -1584 4790
rect -1178 4392 -1118 4790
rect -728 4786 -722 4846
rect -662 4786 -656 4846
rect 1070 4786 1076 4846
rect 1136 4786 1142 4846
rect 1532 4794 1538 4854
rect 1598 4794 1604 4854
rect -722 4392 -662 4786
rect -3928 4332 -662 4392
rect -3926 3910 -3866 4332
rect -3464 3916 -3404 4332
rect -3464 3850 -3404 3856
rect -3010 3910 -2950 4332
rect -2548 3916 -2488 4332
rect -2548 3850 -2488 3856
rect -2094 3916 -2034 4332
rect -2094 3850 -2034 3856
rect -1644 3916 -1584 4332
rect -1644 3850 -1584 3856
rect -1178 3910 -1118 4332
rect -722 3916 -662 4332
rect -488 4724 -428 4730
rect -488 4386 -428 4664
rect 1076 4386 1136 4786
rect 1538 4386 1598 4794
rect 1986 4788 1992 4848
rect 2052 4788 2058 4848
rect 2448 4788 2454 4848
rect 2514 4788 2520 4848
rect 2902 4788 2908 4848
rect 2968 4788 2974 4848
rect 3352 4794 3358 4854
rect 3418 4794 3424 4854
rect 1992 4386 2052 4788
rect 2454 4386 2514 4788
rect 2908 4386 2968 4788
rect 3358 4386 3418 4794
rect 3818 4788 3824 4848
rect 3884 4788 3890 4848
rect 4274 4788 4280 4848
rect 4340 4788 4346 4848
rect 3824 4386 3884 4788
rect 4280 4386 4340 4788
rect 4506 4658 4512 4718
rect 4572 4658 4578 4718
rect -488 4326 4340 4386
rect -488 4044 -428 4326
rect -494 3984 -488 4044
rect -428 3984 -422 4044
rect -722 3850 -662 3856
rect 1076 3916 1136 4326
rect 1076 3850 1136 3856
rect 1538 3914 1598 4326
rect -3926 3844 -3866 3850
rect -3010 3844 -2950 3850
rect -1178 3844 -1118 3850
rect 1538 3848 1598 3854
rect 1992 3914 2052 4326
rect 1992 3848 2052 3854
rect 2454 3914 2514 4326
rect 2454 3848 2514 3854
rect 2908 3914 2968 4326
rect 3358 3920 3418 4326
rect 3358 3854 3418 3860
rect 3824 3916 3884 4326
rect 2908 3848 2968 3854
rect 3824 3850 3884 3856
rect 4280 3916 4340 4326
rect 4512 4382 4572 4658
rect 4512 4322 5598 4382
rect 4512 4056 4572 4322
rect 5498 4193 5598 4322
rect 5494 4103 5503 4193
rect 5593 4103 5602 4193
rect 5498 4098 5598 4103
rect 4512 3990 4572 3996
rect 4280 3850 4340 3856
rect -4680 2448 5090 2476
rect -4680 2362 -4630 2448
rect -4534 2362 -4050 2448
rect -3954 2362 -3450 2448
rect -3354 2362 -2850 2448
rect -2754 2362 -2250 2448
rect -2154 2362 -1650 2448
rect -1554 2362 -1050 2448
rect -954 2362 -450 2448
rect -354 2362 150 2448
rect 246 2362 750 2448
rect 846 2362 1350 2448
rect 1446 2362 1950 2448
rect 2046 2362 2550 2448
rect 2646 2362 3150 2448
rect 3246 2362 3750 2448
rect 3846 2362 4350 2448
rect 4446 2362 4950 2448
rect 5046 2362 5090 2448
rect -4680 2332 5090 2362
rect -4916 2184 -4316 2194
rect -4916 1874 -4316 1884
rect 4716 2184 5316 2194
rect 4716 1874 5316 1884
<< via2 >>
rect -4916 9916 -4316 10216
rect 4716 9916 5316 10216
rect -4064 9656 -3968 9742
rect -3464 9656 -3368 9742
rect -2864 9656 -2768 9742
rect -2264 9656 -2168 9742
rect -1664 9656 -1568 9742
rect -1064 9656 -968 9742
rect -464 9656 -368 9742
rect 136 9656 232 9742
rect 736 9656 832 9742
rect 1336 9656 1432 9742
rect 1936 9656 2032 9742
rect 2536 9656 2632 9742
rect 3136 9656 3232 9742
rect 3736 9656 3832 9742
rect 4156 9656 4252 9742
rect 5503 4103 5593 4193
rect -4630 2362 -4534 2448
rect -4050 2362 -3954 2448
rect -3450 2362 -3354 2448
rect -2850 2362 -2754 2448
rect -2250 2362 -2154 2448
rect -1650 2362 -1554 2448
rect -1050 2362 -954 2448
rect -450 2362 -354 2448
rect 150 2362 246 2448
rect 750 2362 846 2448
rect 1350 2362 1446 2448
rect 1950 2362 2046 2448
rect 2550 2362 2646 2448
rect 3150 2362 3246 2448
rect 3750 2362 3846 2448
rect 4350 2362 4446 2448
rect 4950 2362 5046 2448
rect -4916 1884 -4316 2184
rect 4716 1884 5316 2184
<< metal3 >>
rect -4926 10216 -4306 10221
rect -4926 9916 -4916 10216
rect -4316 9916 -4306 10216
rect -4926 9911 -4306 9916
rect 4706 10216 5326 10221
rect 4706 9916 4716 10216
rect 5316 9916 5326 10216
rect 4706 9911 5326 9916
rect -4078 9742 4278 9756
rect -4078 9656 -4064 9742
rect -3968 9656 -3464 9742
rect -3368 9656 -2864 9742
rect -2768 9656 -2264 9742
rect -2168 9656 -1664 9742
rect -1568 9656 -1064 9742
rect -968 9656 -464 9742
rect -368 9656 136 9742
rect 232 9656 736 9742
rect 832 9656 1336 9742
rect 1432 9656 1936 9742
rect 2032 9656 2536 9742
rect 2632 9656 3136 9742
rect 3232 9656 3736 9742
rect 3832 9656 4156 9742
rect 4252 9656 4278 9742
rect -4078 9646 4278 9656
rect 5498 4197 5598 4198
rect 5493 4099 5499 4197
rect 5597 4099 5603 4197
rect 5498 4098 5598 4099
rect -4680 2448 5090 2476
rect -4680 2362 -4630 2448
rect -4534 2362 -4050 2448
rect -3954 2362 -3450 2448
rect -3354 2362 -2850 2448
rect -2754 2362 -2250 2448
rect -2154 2362 -1650 2448
rect -1554 2362 -1050 2448
rect -954 2362 -450 2448
rect -354 2362 150 2448
rect 246 2362 750 2448
rect 846 2362 1350 2448
rect 1446 2362 1950 2448
rect 2046 2362 2550 2448
rect 2646 2362 3150 2448
rect 3246 2362 3750 2448
rect 3846 2362 4350 2448
rect 4446 2362 4950 2448
rect 5046 2362 5090 2448
rect -4680 2332 5090 2362
rect -4926 2184 -4306 2189
rect -4926 1884 -4916 2184
rect -4316 1884 -4306 2184
rect -4926 1879 -4306 1884
rect 4706 2184 5326 2189
rect 4706 1884 4716 2184
rect 5316 1884 5326 2184
rect 5698 2064 9326 5518
rect 4706 1879 5326 1884
<< via3 >>
rect -4916 9916 -4316 10216
rect 4716 9916 5316 10216
rect -4064 9656 -3968 9742
rect -3464 9656 -3368 9742
rect -2864 9656 -2768 9742
rect -2264 9656 -2168 9742
rect -1664 9656 -1568 9742
rect -1064 9656 -968 9742
rect -464 9656 -368 9742
rect 136 9656 232 9742
rect 736 9656 832 9742
rect 1336 9656 1432 9742
rect 1936 9656 2032 9742
rect 2536 9656 2632 9742
rect 3136 9656 3232 9742
rect 3736 9656 3832 9742
rect 4156 9656 4252 9742
rect 5499 4193 5597 4197
rect 5499 4103 5503 4193
rect 5503 4103 5593 4193
rect 5593 4103 5597 4193
rect 5499 4099 5597 4103
rect -4630 2362 -4534 2448
rect -4050 2362 -3954 2448
rect -3450 2362 -3354 2448
rect -2850 2362 -2754 2448
rect -2250 2362 -2154 2448
rect -1650 2362 -1554 2448
rect -1050 2362 -954 2448
rect -450 2362 -354 2448
rect 150 2362 246 2448
rect 750 2362 846 2448
rect 1350 2362 1446 2448
rect 1950 2362 2046 2448
rect 2550 2362 2646 2448
rect 3150 2362 3246 2448
rect 3750 2362 3846 2448
rect 4350 2362 4446 2448
rect 4950 2362 5046 2448
rect -4916 1884 -4316 2184
rect 4716 1884 5316 2184
<< metal4 >>
rect -5100 10216 9448 10400
rect -5100 9916 -4916 10216
rect -4316 9916 4716 10216
rect 5316 9916 9448 10216
rect -5100 9742 9448 9916
rect -5100 9656 -4064 9742
rect -3968 9656 -3464 9742
rect -3368 9656 -2864 9742
rect -2768 9656 -2264 9742
rect -2168 9656 -1664 9742
rect -1568 9656 -1064 9742
rect -968 9656 -464 9742
rect -368 9656 136 9742
rect 232 9656 736 9742
rect 832 9656 1336 9742
rect 1432 9656 1936 9742
rect 2032 9656 2536 9742
rect 2632 9656 3136 9742
rect 3232 9656 3736 9742
rect 3832 9656 4156 9742
rect 4252 9656 9448 9742
rect -5100 9600 9448 9656
rect 5974 5144 9288 5244
rect 5974 4554 6074 5144
rect 6310 4554 6410 5144
rect 5974 4454 6410 4554
rect 5974 4340 6074 4454
rect 6310 4340 6410 4454
rect 6688 4790 8232 4890
rect 6688 4198 6788 4790
rect 7408 4198 7508 4790
rect 8130 4198 8231 4790
rect 8476 4555 8578 5144
rect 8478 4550 8578 4555
rect 8850 4550 8950 5144
rect 9188 5089 9288 5144
rect 9188 4594 9291 5089
rect 9188 4550 9288 4594
rect 8478 4450 9288 4550
rect 8478 4300 8578 4450
rect 8850 4338 8950 4450
rect 9188 4300 9288 4450
rect 5498 4197 9450 4198
rect 5498 4099 5499 4197
rect 5597 4099 9450 4197
rect 5498 4098 9450 4099
rect 5974 3852 6074 3962
rect 6310 3852 6410 3962
rect 5974 3752 6410 3852
rect 5974 3146 6074 3752
rect 6310 3146 6410 3752
rect 5974 3046 6410 3146
rect 5974 2500 6074 3046
rect 6310 2500 6410 3046
rect 6688 3496 6788 4098
rect 7408 3496 7508 4098
rect 8130 3496 8231 4098
rect 6688 3396 8231 3496
rect 6688 2796 6788 3396
rect 7408 2796 7508 3396
rect 8130 2796 8231 3396
rect 8478 3846 8578 4000
rect 8850 3846 8950 3962
rect 9188 3846 9288 4000
rect 8478 3746 9288 3846
rect 8478 3154 8578 3746
rect 8850 3154 8950 3746
rect 9188 3154 9288 3746
rect 8478 3054 9288 3154
rect 8478 2995 8578 3054
rect 6688 2696 8232 2796
rect 8476 2500 8578 2995
rect 8850 2500 8950 3054
rect 9188 3035 9288 3054
rect 9188 2500 9291 3035
rect -5100 2448 9448 2500
rect -5100 2362 -4630 2448
rect -4534 2362 -4050 2448
rect -3954 2362 -3450 2448
rect -3354 2362 -2850 2448
rect -2754 2362 -2250 2448
rect -2154 2362 -1650 2448
rect -1554 2362 -1050 2448
rect -954 2362 -450 2448
rect -354 2362 150 2448
rect 246 2362 750 2448
rect 846 2362 1350 2448
rect 1446 2362 1950 2448
rect 2046 2362 2550 2448
rect 2646 2362 3150 2448
rect 3246 2362 3750 2448
rect 3846 2362 4350 2448
rect 4446 2362 4950 2448
rect 5046 2362 9448 2448
rect -5100 2184 9448 2362
rect -5100 1884 -4916 2184
rect -4316 1884 4716 2184
rect 5316 1884 9448 2184
rect -5100 1700 9448 1884
rect 8478 1696 8578 1700
use sky130_fd_pr__cap_mim_m3_1_FAR8MD  sky130_fd_pr__cap_mim_m3_1_FAR8MD_0
timestamp 1623971255
transform 1 0 7508 0 1 3800
box -1788 -1700 1787 1700
use sky130_fd_pr__pfet_01v8_hvt_8Q5PU3  sky130_fd_pr__pfet_01v8_hvt_8Q5PU3_0
timestamp 1623971255
transform 1 0 -2288 0 1 5605
box -2355 -700 2355 700
use sky130_fd_pr__pfet_01v8_hvt_8Q5PU3  sky130_fd_pr__pfet_01v8_hvt_8Q5PU3_1
timestamp 1623971255
transform 1 0 2712 0 1 5605
box -2355 -700 2355 700
use sky130_fd_pr__pfet_01v8_hvt_GK2P2M  sky130_fd_pr__pfet_01v8_hvt_GK2P2M_0
timestamp 1623971255
transform 1 0 103 0 1 8070
box -4187 -900 4187 900
use sky130_fd_pr__nfet_01v8_V6PJ6N  sky130_fd_pr__nfet_01v8_V6PJ6N_2
timestamp 1623971255
transform 1 0 2711 0 1 3612
box -2319 -188 2319 188
use sky130_fd_pr__nfet_01v8_V6PJ6N  sky130_fd_pr__nfet_01v8_V6PJ6N_1
timestamp 1623971255
transform 1 0 -2289 0 1 3612
box -2319 -188 2319 188
use sky130_fd_pr__nfet_01v8_V6PJ6N  sky130_fd_pr__nfet_01v8_V6PJ6N_0
timestamp 1623971255
transform 1 0 -2289 0 1 2944
box -2319 -188 2319 188
<< labels >>
flabel metal4 -2300 2102 -2280 2122 1 FreeSans 480 0 0 0 VSS
flabel metal4 -2534 10006 -2500 10030 1 FreeSans 480 0 0 0 VDD
flabel metal2 -3700 4356 -3686 4370 1 FreeSans 480 0 0 0 vin
flabel metal1 -3698 2662 -3690 2672 1 FreeSans 480 0 0 0 vbiasn
flabel metal2 -3228 7078 -3218 7084 1 FreeSans 480 0 0 0 vbiasp
flabel metal2 4126 4350 4138 4364 1 FreeSans 480 0 0 0 voutcs
flabel metal2 4532 4380 4544 4390 1 FreeSans 480 0 0 0 vout
flabel metal1 -4134 3252 -4122 3270 1 FreeSans 480 0 0 0 csinvn
flabel metal2 -3584 6480 -3574 6494 1 FreeSans 480 0 0 0 csinvp
<< properties >>
string FIXED_BBOX -4972 1328 5372 4032
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nwell >>
rect -968 -300 968 300
<< pmos >>
rect -874 -200 -674 200
rect -616 -200 -416 200
rect -358 -200 -158 200
rect -100 -200 100 200
rect 158 -200 358 200
rect 416 -200 616 200
rect 674 -200 874 200
<< pdiff >>
rect -932 188 -874 200
rect -932 -188 -920 188
rect -886 -188 -874 188
rect -932 -200 -874 -188
rect -674 188 -616 200
rect -674 -188 -662 188
rect -628 -188 -616 188
rect -674 -200 -616 -188
rect -416 188 -358 200
rect -416 -188 -404 188
rect -370 -188 -358 188
rect -416 -200 -358 -188
rect -158 188 -100 200
rect -158 -188 -146 188
rect -112 -188 -100 188
rect -158 -200 -100 -188
rect 100 188 158 200
rect 100 -188 112 188
rect 146 -188 158 188
rect 100 -200 158 -188
rect 358 188 416 200
rect 358 -188 370 188
rect 404 -188 416 188
rect 358 -200 416 -188
rect 616 188 674 200
rect 616 -188 628 188
rect 662 -188 674 188
rect 616 -200 674 -188
rect 874 188 932 200
rect 874 -188 886 188
rect 920 -188 932 188
rect 874 -200 932 -188
<< pdiffc >>
rect -920 -188 -886 188
rect -662 -188 -628 188
rect -404 -188 -370 188
rect -146 -188 -112 188
rect 112 -188 146 188
rect 370 -188 404 188
rect 628 -188 662 188
rect 886 -188 920 188
<< poly >>
rect -840 281 -708 297
rect -840 264 -824 281
rect -874 247 -824 264
rect -724 264 -708 281
rect -582 281 -450 297
rect -582 264 -566 281
rect -724 247 -674 264
rect -874 200 -674 247
rect -616 247 -566 264
rect -466 264 -450 281
rect -324 281 -192 297
rect -324 264 -308 281
rect -466 247 -416 264
rect -616 200 -416 247
rect -358 247 -308 264
rect -208 264 -192 281
rect -66 281 66 297
rect -66 264 -50 281
rect -208 247 -158 264
rect -358 200 -158 247
rect -100 247 -50 264
rect 50 264 66 281
rect 192 281 324 297
rect 192 264 208 281
rect 50 247 100 264
rect -100 200 100 247
rect 158 247 208 264
rect 308 264 324 281
rect 450 281 582 297
rect 450 264 466 281
rect 308 247 358 264
rect 158 200 358 247
rect 416 247 466 264
rect 566 264 582 281
rect 708 281 840 297
rect 708 264 724 281
rect 566 247 616 264
rect 416 200 616 247
rect 674 247 724 264
rect 824 264 840 281
rect 824 247 874 264
rect 674 200 874 247
rect -874 -247 -674 -200
rect -874 -264 -824 -247
rect -840 -281 -824 -264
rect -724 -264 -674 -247
rect -616 -247 -416 -200
rect -616 -264 -566 -247
rect -724 -281 -708 -264
rect -840 -297 -708 -281
rect -582 -281 -566 -264
rect -466 -264 -416 -247
rect -358 -247 -158 -200
rect -358 -264 -308 -247
rect -466 -281 -450 -264
rect -582 -297 -450 -281
rect -324 -281 -308 -264
rect -208 -264 -158 -247
rect -100 -247 100 -200
rect -100 -264 -50 -247
rect -208 -281 -192 -264
rect -324 -297 -192 -281
rect -66 -281 -50 -264
rect 50 -264 100 -247
rect 158 -247 358 -200
rect 158 -264 208 -247
rect 50 -281 66 -264
rect -66 -297 66 -281
rect 192 -281 208 -264
rect 308 -264 358 -247
rect 416 -247 616 -200
rect 416 -264 466 -247
rect 308 -281 324 -264
rect 192 -297 324 -281
rect 450 -281 466 -264
rect 566 -264 616 -247
rect 674 -247 874 -200
rect 674 -264 724 -247
rect 566 -281 582 -264
rect 450 -297 582 -281
rect 708 -281 724 -264
rect 824 -264 874 -247
rect 824 -281 840 -264
rect 708 -297 840 -281
<< polycont >>
rect -824 247 -724 281
rect -566 247 -466 281
rect -308 247 -208 281
rect -50 247 50 281
rect 208 247 308 281
rect 466 247 566 281
rect 724 247 824 281
rect -824 -281 -724 -247
rect -566 -281 -466 -247
rect -308 -281 -208 -247
rect -50 -281 50 -247
rect 208 -281 308 -247
rect 466 -281 566 -247
rect 724 -281 824 -247
<< locali >>
rect -840 247 -824 281
rect -724 247 -708 281
rect -582 247 -566 281
rect -466 247 -450 281
rect -324 247 -308 281
rect -208 247 -192 281
rect -66 247 -50 281
rect 50 247 66 281
rect 192 247 208 281
rect 308 247 324 281
rect 450 247 466 281
rect 566 247 582 281
rect 708 247 724 281
rect 824 247 840 281
rect -920 188 -886 204
rect -920 -204 -886 -188
rect -662 188 -628 204
rect -662 -204 -628 -188
rect -404 188 -370 204
rect -404 -204 -370 -188
rect -146 188 -112 204
rect -146 -204 -112 -188
rect 112 188 146 204
rect 112 -204 146 -188
rect 370 188 404 204
rect 370 -204 404 -188
rect 628 188 662 204
rect 628 -204 662 -188
rect 886 188 920 204
rect 886 -204 920 -188
rect -840 -281 -824 -247
rect -724 -281 -708 -247
rect -582 -281 -566 -247
rect -466 -281 -450 -247
rect -324 -281 -308 -247
rect -208 -281 -192 -247
rect -66 -281 -50 -247
rect 50 -281 66 -247
rect 192 -281 208 -247
rect 308 -281 324 -247
rect 450 -281 466 -247
rect 566 -281 582 -247
rect 708 -281 724 -247
rect 824 -281 840 -247
<< viali >>
rect -816 247 -732 281
rect -558 247 -474 281
rect -300 247 -216 281
rect -42 247 42 281
rect 216 247 300 281
rect 474 247 558 281
rect 732 247 816 281
rect -920 -188 -886 188
rect -662 -188 -628 188
rect -404 -188 -370 188
rect -146 -188 -112 188
rect 112 -188 146 188
rect 370 -188 404 188
rect 628 -188 662 188
rect 886 -188 920 188
rect -816 -281 -732 -247
rect -558 -281 -474 -247
rect -300 -281 -216 -247
rect -42 -281 42 -247
rect 216 -281 300 -247
rect 474 -281 558 -247
rect 732 -281 816 -247
<< metal1 >>
rect -828 281 -720 287
rect -828 247 -816 281
rect -732 247 -720 281
rect -828 241 -720 247
rect -570 281 -462 287
rect -570 247 -558 281
rect -474 247 -462 281
rect -570 241 -462 247
rect -312 281 -204 287
rect -312 247 -300 281
rect -216 247 -204 281
rect -312 241 -204 247
rect -54 281 54 287
rect -54 247 -42 281
rect 42 247 54 281
rect -54 241 54 247
rect 204 281 312 287
rect 204 247 216 281
rect 300 247 312 281
rect 204 241 312 247
rect 462 281 570 287
rect 462 247 474 281
rect 558 247 570 281
rect 462 241 570 247
rect 720 281 828 287
rect 720 247 732 281
rect 816 247 828 281
rect 720 241 828 247
rect -926 188 -880 200
rect -926 -188 -920 188
rect -886 -188 -880 188
rect -926 -200 -880 -188
rect -668 188 -622 200
rect -668 -188 -662 188
rect -628 -188 -622 188
rect -668 -200 -622 -188
rect -410 188 -364 200
rect -410 -188 -404 188
rect -370 -188 -364 188
rect -410 -200 -364 -188
rect -152 188 -106 200
rect -152 -188 -146 188
rect -112 -188 -106 188
rect -152 -200 -106 -188
rect 106 188 152 200
rect 106 -188 112 188
rect 146 -188 152 188
rect 106 -200 152 -188
rect 364 188 410 200
rect 364 -188 370 188
rect 404 -188 410 188
rect 364 -200 410 -188
rect 622 188 668 200
rect 622 -188 628 188
rect 662 -188 668 188
rect 622 -200 668 -188
rect 880 188 926 200
rect 880 -188 886 188
rect 920 -188 926 188
rect 880 -200 926 -188
rect -828 -247 -720 -241
rect -828 -281 -816 -247
rect -732 -281 -720 -247
rect -828 -287 -720 -281
rect -570 -247 -462 -241
rect -570 -281 -558 -247
rect -474 -281 -462 -247
rect -570 -287 -462 -281
rect -312 -247 -204 -241
rect -312 -281 -300 -247
rect -216 -281 -204 -247
rect -312 -287 -204 -281
rect -54 -247 54 -241
rect -54 -281 -42 -247
rect 42 -281 54 -247
rect -54 -287 54 -281
rect 204 -247 312 -241
rect 204 -281 216 -247
rect 300 -281 312 -247
rect 204 -287 312 -281
rect 462 -247 570 -241
rect 462 -281 474 -247
rect 558 -281 570 -247
rect 462 -287 570 -281
rect 720 -247 828 -241
rect 720 -281 732 -247
rect 816 -281 828 -247
rect 720 -287 828 -281
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string parameters w 2 l 1 m 1 nf 7 diffcov 100 polycov 60 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1624136344
<< nwell >>
rect -12082 15478 -10232 16318
rect -8617 15502 -7946 15800
rect -8617 15479 -8084 15502
rect -7962 15479 -7946 15502
<< pwell >>
rect -8558 15406 -8084 15421
rect -11841 14764 -10108 15384
rect -8558 15239 -7981 15406
<< viali >>
rect -8052 15430 -8004 15478
rect -7950 15434 -7902 15482
<< metal1 >>
rect 47792 27680 48000 27710
rect -1414 27642 -1354 27648
rect -1414 16408 -1354 27582
rect 47792 27564 47824 27680
rect 47022 25478 47376 25538
rect 47792 25514 48000 27564
rect 48306 27680 48488 27710
rect 48462 27564 48488 27680
rect 48306 25497 48488 27564
rect 47022 23538 47082 25478
rect 47244 23874 47250 23934
rect 47310 23874 47316 23934
rect 47022 23478 47802 23538
rect 48682 23478 50478 23538
rect 46972 21860 46978 21920
rect 47038 21860 47310 21920
rect -11720 16348 -10286 16408
rect -9282 16348 -8730 16408
rect -8670 16348 -8664 16408
rect -1420 16348 -1414 16408
rect -1354 16348 -1348 16408
rect -8340 15714 -8100 15810
rect -13304 15478 -13204 15484
rect -8299 15478 -7992 15484
rect -13204 15402 -12676 15462
rect -8299 15430 -8052 15478
rect -8004 15430 -7992 15478
rect -8299 15424 -7992 15430
rect -7962 15482 -7734 15488
rect -7962 15434 -7950 15482
rect -7902 15434 -7734 15482
rect -7962 15428 -7734 15434
rect -12742 15382 -12732 15402
rect -10142 15380 -10130 15400
rect -13304 15372 -13204 15378
rect -12478 14976 -12418 15256
rect -12478 14910 -12418 14916
rect -9878 14944 -9818 15278
rect -8340 15170 -8100 15266
rect -9878 14878 -9818 14884
rect -10012 14777 -10006 14837
rect -9946 14777 -9748 14837
rect -10508 14712 -10502 14730
rect -1792 14712 -1732 14718
rect -11698 14652 -10086 14712
rect -9152 14652 -8724 14712
rect -8664 14652 -8658 14712
rect -1732 14652 -1294 14712
rect -1792 14646 -1732 14652
rect 48494 8574 48554 8578
rect 48494 8514 49142 8574
rect 50076 8546 50476 23478
rect 50938 9088 50944 9148
rect 51004 9088 51010 9148
rect 48358 7491 48364 7551
rect 48424 7491 48430 7551
rect 48364 6090 48424 7491
rect 48494 6610 48554 8514
rect 50944 7650 51004 9088
rect 50812 7590 51004 7650
rect 49766 6818 52704 6878
rect 48494 6550 48854 6610
rect 48358 6030 48364 6090
rect 48424 6030 48430 6090
rect 8274 5144 8280 5204
rect 8340 5144 8346 5204
rect 3944 4926 4244 4986
rect 8280 4788 8340 5144
rect 48494 4610 48554 6550
rect 50810 5626 51006 5686
rect 57932 4926 58226 4986
rect 49930 4854 52710 4914
rect 48494 4550 48994 4610
rect 48494 2520 48554 4550
rect 49960 2854 52704 2914
rect 48494 2462 49148 2520
rect 48498 2460 49148 2462
rect 50008 764 52706 824
<< via1 >>
rect -1414 27582 -1354 27642
rect 47824 27564 48000 27680
rect 48306 27564 48462 27680
rect 47250 23874 47310 23934
rect 46978 21860 47038 21920
rect -8730 16348 -8670 16408
rect -1414 16348 -1354 16408
rect -13304 15378 -13204 15478
rect -12478 14916 -12418 14976
rect -9878 14884 -9818 14944
rect -10006 14777 -9946 14837
rect -8724 14652 -8664 14712
rect -1792 14652 -1732 14712
rect 50944 9088 51004 9148
rect 48364 7491 48424 7551
rect 48364 6030 48424 6090
rect 8280 5144 8340 5204
<< metal2 >>
rect 47796 27680 48490 27702
rect -1414 27642 -1354 27651
rect -1420 27582 -1414 27642
rect -1354 27582 -1348 27642
rect -1414 27573 -1354 27582
rect 47796 27564 47824 27680
rect 48462 27564 48490 27680
rect 47796 27536 48490 27564
rect 48230 24604 48398 24664
rect 48458 24604 48467 24664
rect 47615 24455 47624 24515
rect 47684 24455 47782 24515
rect 47250 23934 47310 23940
rect 42831 23874 42840 23934
rect 42900 23874 47250 23934
rect 47250 23868 47310 23874
rect 47867 22604 47876 22664
rect 47936 22604 48046 22664
rect 48514 22455 48656 22515
rect 48716 22455 48725 22515
rect 49519 22328 49579 24074
rect 46978 21920 47038 21926
rect 42815 21860 42824 21920
rect 42884 21860 46978 21920
rect 46978 21854 47038 21860
rect 40179 21696 40269 21700
rect 36254 21691 40274 21696
rect 36254 21601 40179 21691
rect 40269 21601 40274 21691
rect 36254 21596 40274 21601
rect 11206 18913 11306 18918
rect 11202 18823 11211 18913
rect 11301 18823 11310 18913
rect -8730 16408 -8670 16414
rect -1414 16408 -1354 16414
rect -8670 16348 -1414 16408
rect -8730 16342 -8670 16348
rect -1414 16342 -1354 16348
rect 10953 16318 10962 16418
rect 11062 16318 11071 16418
rect -13299 15478 -13209 15482
rect -13310 15378 -13304 15478
rect -13204 15378 -13198 15478
rect -13299 15374 -13209 15378
rect -10629 15325 -10620 15385
rect -10560 15325 -10006 15385
rect -1933 15226 -1924 15286
rect -1864 15226 -1855 15286
rect -12484 14916 -12478 14976
rect -12418 14916 -12412 14976
rect -13467 14610 -13377 14614
rect -12478 14610 -12418 14916
rect -9884 14884 -9878 14944
rect -9818 14884 -9812 14944
rect -10006 14837 -9946 14843
rect -10838 14777 -10006 14837
rect -10006 14771 -9946 14777
rect -13472 14605 -12418 14610
rect -13472 14515 -13467 14605
rect -13377 14515 -12418 14605
rect -13472 14510 -12418 14515
rect -13467 14506 -13377 14510
rect -9878 13016 -9818 14884
rect -1924 14838 -1864 15226
rect 10962 15101 11062 16318
rect 11206 15882 11306 18823
rect 36254 16193 36354 21596
rect 40179 21592 40269 21596
rect 65088 18913 65188 18918
rect 65084 18823 65093 18913
rect 65183 18823 65192 18913
rect 36250 16103 36259 16193
rect 36349 16103 36358 16193
rect 36254 16098 36354 16103
rect 11197 15782 11206 15882
rect 11306 15782 11315 15882
rect 10958 15011 10967 15101
rect 11057 15011 11066 15101
rect 10962 15006 11062 15011
rect -8360 14778 -1864 14838
rect 11206 14812 11306 15782
rect -8724 14712 -8664 14718
rect 11197 14712 11206 14812
rect 11306 14712 11315 14812
rect 65088 14738 65188 18823
rect -8664 14652 -1792 14712
rect -1732 14652 -1726 14712
rect -8724 14646 -8664 14652
rect 65079 14638 65088 14738
rect 65188 14638 65197 14738
rect 36456 13712 36556 13721
rect 39253 13712 39343 13716
rect 36556 13707 39348 13712
rect 36556 13617 39253 13707
rect 39343 13617 39348 13707
rect 36556 13612 39348 13617
rect 36456 13603 36556 13612
rect 39253 13608 39343 13612
rect -9878 12947 -9818 12956
rect 36060 9390 36160 9399
rect 39009 9390 39099 9394
rect 36056 9290 36060 9390
rect 36160 9385 39104 9390
rect 36160 9295 39009 9385
rect 39099 9295 39104 9385
rect 36160 9290 39104 9295
rect 36060 9281 36160 9290
rect 39009 9286 39099 9290
rect 35833 9172 35935 9176
rect 35828 9167 51026 9172
rect 35828 9065 35833 9167
rect 35935 9148 51026 9167
rect 35935 9088 50944 9148
rect 51004 9088 51026 9148
rect 35935 9065 51026 9088
rect 35828 9060 51026 9065
rect 35833 9056 35935 9060
rect 49704 7640 49822 7700
rect 49882 7640 49891 7700
rect 48364 7551 48424 7557
rect 48424 7491 49184 7551
rect 48364 7485 48424 7491
rect 11382 7198 11442 7207
rect 9888 7138 11382 7198
rect 62341 7138 62350 7198
rect 62410 7138 62660 7198
rect 11382 7129 11442 7138
rect 50834 6944 51160 7004
rect 46253 6112 46343 6116
rect 46248 6107 48434 6112
rect 46248 6017 46253 6107
rect 46343 6090 48434 6107
rect 46343 6030 48364 6090
rect 48424 6030 48434 6090
rect 46343 6017 48434 6030
rect 46248 6012 48434 6017
rect 46253 6008 46343 6012
rect 49297 5676 49306 5736
rect 49366 5676 49510 5736
rect 49931 5527 49940 5587
rect 50000 5527 50009 5587
rect 8280 5204 8340 5210
rect 8271 5144 8280 5204
rect 8340 5144 8349 5204
rect 8280 5138 8340 5144
rect 49293 3676 49302 3736
rect 49362 3676 49472 3736
rect 49940 3527 50082 3587
rect 50142 3527 50151 3587
rect 50945 3400 51005 5146
rect 46279 1708 46288 1768
rect 46348 1708 46357 1768
rect 8042 1566 9100 1626
rect 8042 582 8102 1566
rect 46288 1497 46348 1708
rect 49734 1586 49828 1646
rect 49888 1586 49897 1646
rect 51100 1596 51160 6944
rect 66017 4876 66026 4936
rect 66086 4876 66095 4936
rect 66026 3818 66086 4876
rect 65964 3758 66086 3818
rect 62153 2933 62243 2942
rect 62243 2860 62414 2920
rect 62153 2834 62243 2843
rect 50940 1536 51160 1596
rect 46288 1437 49196 1497
rect 8033 522 8042 582
rect 8102 522 8111 582
<< via2 >>
rect -1414 27582 -1354 27642
rect 47824 27564 48000 27680
rect 48000 27564 48306 27680
rect 48306 27564 48462 27680
rect 48398 24604 48458 24664
rect 47624 24455 47684 24515
rect 42840 23874 42900 23934
rect 47876 22604 47936 22664
rect 48656 22455 48716 22515
rect 42824 21860 42884 21920
rect 40179 21601 40269 21691
rect 11211 18823 11301 18913
rect 10962 16318 11062 16418
rect -13299 15383 -13209 15473
rect -10620 15325 -10560 15385
rect -1924 15226 -1864 15286
rect -13467 14515 -13377 14605
rect 65093 18823 65183 18913
rect 36259 16103 36349 16193
rect 11206 15782 11306 15882
rect 10967 15011 11057 15101
rect 11206 14712 11306 14812
rect 65088 14638 65188 14738
rect 36456 13612 36556 13712
rect 39253 13617 39343 13707
rect -9878 12956 -9818 13016
rect 36060 9290 36160 9390
rect 39009 9295 39099 9385
rect 35833 9065 35935 9167
rect 49822 7640 49882 7700
rect 11382 7138 11442 7198
rect 62350 7138 62410 7198
rect 46253 6017 46343 6107
rect 49306 5676 49366 5736
rect 49940 5527 50000 5587
rect 8280 5144 8340 5204
rect 49302 3676 49362 3736
rect 50082 3527 50142 3587
rect 46288 1708 46348 1768
rect 49828 1586 49888 1646
rect 66026 4876 66086 4936
rect 62153 2843 62243 2933
rect 8042 522 8102 582
<< metal3 >>
rect 47796 27680 48490 27702
rect -1436 27647 -1330 27668
rect -1436 27583 -1419 27647
rect -1349 27583 -1330 27647
rect -1436 27582 -1414 27583
rect -1354 27582 -1330 27583
rect -1436 27562 -1330 27582
rect 47796 27564 47824 27680
rect 48462 27564 48490 27680
rect 47796 27536 48490 27564
rect 38288 27302 38888 27308
rect 37303 26378 38288 26434
rect 41068 27302 41668 27308
rect 38888 26378 41068 26434
rect 41668 26378 42904 26434
rect 37303 25834 42904 26378
rect 37303 25000 37903 25834
rect 36728 24400 36734 25000
rect 37334 24400 37903 25000
rect 36468 23705 36568 23706
rect 36463 23607 36469 23705
rect 36567 23607 36573 23705
rect 36468 20168 36568 23607
rect 37303 22924 37903 24400
rect 39700 23708 39800 23958
rect 39508 23705 39608 23706
rect 39503 23607 39509 23705
rect 39607 23607 39613 23705
rect 39700 23608 40274 23708
rect 40402 23706 40502 23944
rect 42304 23939 42904 25834
rect 43504 24440 43510 25040
rect 48378 24664 51894 24688
rect 48378 24604 48398 24664
rect 48458 24604 51894 24664
rect 48378 24588 51894 24604
rect 46576 24534 46676 24540
rect 46676 24515 47704 24534
rect 46676 24455 47624 24515
rect 47684 24455 47704 24515
rect 46676 24434 47704 24455
rect 46576 24428 46676 24434
rect 42304 23934 42905 23939
rect 42304 23874 42840 23934
rect 42900 23874 42905 23934
rect 42304 23869 42905 23874
rect 41563 23712 41661 23717
rect 42094 23712 42194 23718
rect 41562 23711 42094 23712
rect 39508 23306 39608 23607
rect 36732 22324 36738 22924
rect 37338 22324 37903 22924
rect 37270 22322 37903 22324
rect 37303 21496 37903 22322
rect 40174 21691 40274 23608
rect 40396 23606 40402 23706
rect 40502 23606 40508 23706
rect 41562 23613 41563 23711
rect 41661 23613 42094 23711
rect 41562 23612 42094 23613
rect 41563 23607 41661 23612
rect 42094 23606 42194 23612
rect 40174 21601 40179 21691
rect 40269 21601 40274 21691
rect 40174 21596 40274 21601
rect 42304 22912 42904 23869
rect 42304 22312 42914 22912
rect 43514 22312 43520 22912
rect 46402 22664 47952 22684
rect 46402 22604 47876 22664
rect 47936 22604 47952 22664
rect 46402 22584 47952 22604
rect 42304 21920 42904 22312
rect 46402 22156 46502 22584
rect 48640 22515 49860 22532
rect 48640 22455 48656 22515
rect 48716 22455 49860 22515
rect 48640 22432 49860 22455
rect 46402 22046 46504 22156
rect 42304 21860 42824 21920
rect 42884 21860 42904 21920
rect 38277 21496 38879 21498
rect 41047 21496 41649 21498
rect 42304 21496 42904 21860
rect 37303 20896 42904 21496
rect 44725 21200 45327 21206
rect 37304 20593 42896 20896
rect 46404 21103 46504 22046
rect 49760 21700 49860 22432
rect 49760 21594 49860 21600
rect 47028 21132 47628 21138
rect 46399 21005 46405 21103
rect 46503 21005 46509 21103
rect 46404 21004 46504 21005
rect 37304 20589 43176 20593
rect 44152 20589 44258 20593
rect 44725 20589 45327 20598
rect 46654 20589 46804 20590
rect 37304 20584 47028 20589
rect 37297 20532 47028 20584
rect 49808 21132 50408 21138
rect 47628 20532 49808 20588
rect 51794 21066 51894 24588
rect 52138 23614 52144 23714
rect 52244 23614 52250 23714
rect 51788 20966 51794 21066
rect 51894 20966 51900 21066
rect 50408 20532 51393 20588
rect 36468 19829 36572 20168
rect 37297 19984 51393 20532
rect 36467 19731 36473 19829
rect 36571 19731 36577 19829
rect 11036 18913 11638 18918
rect 11036 18823 11211 18913
rect 11301 18823 11638 18913
rect 11036 18818 11638 18823
rect 36468 17152 36572 19731
rect 37297 18950 37897 19984
rect 39072 19730 39078 19830
rect 39178 19730 46764 19830
rect 36710 18350 36716 18950
rect 37316 18350 37897 18950
rect 36468 17048 36852 17152
rect 10957 16418 11067 16423
rect 10957 16318 10962 16418
rect 11062 16318 11067 16418
rect 11464 16322 36558 16422
rect 10957 16313 11067 16318
rect 36254 16193 36354 16198
rect 36254 16103 36259 16193
rect 36349 16103 36354 16193
rect 11201 15882 11311 15887
rect 11201 15782 11206 15882
rect 11306 15782 36158 15882
rect 11201 15777 11311 15782
rect -13304 15473 -13204 15478
rect -13304 15383 -13299 15473
rect -13209 15383 -13204 15473
rect -13304 14732 -13204 15383
rect -10642 15385 -10542 15410
rect -10642 15325 -10620 15385
rect -10560 15325 -10542 15385
rect -10642 14732 -10542 15325
rect -1950 15286 35940 15316
rect -1950 15226 -1924 15286
rect -1864 15226 35940 15286
rect -1950 15204 35940 15226
rect -13304 14632 -10542 14732
rect -2396 15101 11062 15106
rect -2396 15011 10967 15101
rect 11057 15011 11062 15101
rect -2396 15006 11062 15011
rect -13472 14605 -13372 14610
rect -13472 14515 -13467 14605
rect -13377 14515 -13372 14605
rect -13472 10875 -13372 14515
rect -13477 10777 -13471 10875
rect -13373 10777 -13367 10875
rect -13472 10776 -13372 10777
rect -13304 3637 -13204 14632
rect -11340 14342 -10740 14348
rect -12325 13742 -11340 13798
rect -8560 14342 -7960 14348
rect -10740 13742 -8560 13798
rect -6972 14344 -6372 14350
rect -7736 13798 -6972 13800
rect -7960 13744 -6972 13798
rect -4192 14344 -3592 14350
rect -6372 13744 -4192 13800
rect -3592 13744 -2607 13800
rect -7960 13742 -2607 13744
rect -12325 13200 -2607 13742
rect -12325 13198 -7666 13200
rect -13108 13033 -13008 13034
rect -13113 12935 -13107 13033
rect -13009 12935 -13003 13033
rect -13108 12772 -13006 12935
rect -13106 9154 -13006 12772
rect -12325 12164 -11725 13198
rect -10580 12934 -10574 13034
rect -10474 13016 -7214 13034
rect -10474 12956 -9878 13016
rect -9818 12956 -7214 13016
rect -10474 12934 -7214 12956
rect -12912 11564 -12906 12164
rect -12306 11564 -11725 12164
rect -12325 10086 -11725 11564
rect -9964 10878 -9864 12934
rect -7314 12716 -7214 12934
rect -3207 12166 -2607 13200
rect -2396 12904 -2296 15006
rect 11201 14812 11311 14817
rect 10974 14810 11206 14812
rect -1756 14712 11206 14810
rect 11306 14712 11311 14812
rect -1756 14710 11311 14712
rect -2402 12804 -2396 12904
rect -2296 12804 -2290 12904
rect -3207 11566 -2626 12166
rect -2026 11566 -2020 12166
rect -10156 10875 -10056 10876
rect -10161 10777 -10155 10875
rect -10057 10777 -10051 10875
rect -9964 10778 -9390 10878
rect -9262 10876 -9162 11114
rect -8101 10882 -8003 10887
rect -7570 10882 -7470 10888
rect -8102 10881 -7570 10882
rect -10156 10588 -10056 10777
rect -10156 10476 -10002 10588
rect -9490 10492 -9390 10778
rect -9268 10776 -9262 10876
rect -9162 10776 -9156 10876
rect -8102 10783 -8101 10881
rect -8003 10783 -7570 10881
rect -8102 10782 -7570 10783
rect -5764 10878 -5664 11128
rect -5956 10875 -5856 10876
rect -8101 10777 -8003 10782
rect -7570 10776 -7470 10782
rect -5961 10777 -5955 10875
rect -5857 10777 -5851 10875
rect -5764 10778 -5190 10878
rect -5062 10876 -4962 11114
rect -3901 10880 -3803 10885
rect -3370 10880 -3270 10886
rect -3902 10879 -3370 10880
rect -7192 10492 -7190 10684
rect -5956 10476 -5856 10777
rect -5290 10684 -5190 10778
rect -5068 10776 -5062 10876
rect -4962 10776 -4956 10876
rect -3902 10781 -3901 10879
rect -3803 10781 -3370 10879
rect -3902 10780 -3370 10781
rect -3901 10775 -3803 10780
rect -3370 10774 -3270 10780
rect -5290 10492 -5192 10684
rect -12922 9486 -12916 10086
rect -12316 9486 -11725 10086
rect -13106 9054 -12632 9154
rect -13100 8711 -13000 8712
rect -13105 8613 -13099 8711
rect -13001 8613 -12995 8711
rect -13309 3539 -13303 3637
rect -13205 3539 -13199 3637
rect -13304 3538 -13204 3539
rect -13100 1627 -13000 8613
rect -12732 5665 -12632 9054
rect -12325 8460 -11725 9486
rect -10102 8712 -10002 10476
rect -3207 10088 -2607 11566
rect -1756 11018 -1656 14710
rect 11201 14707 11311 14710
rect -3207 9488 -2616 10088
rect -2016 9488 -2010 10088
rect -7192 8712 -7092 9154
rect -10510 8612 -10504 8712
rect -10404 8612 -7092 8712
rect -6953 8462 -6351 8464
rect -4183 8462 -3581 8464
rect -3207 8462 -2607 9488
rect -1758 8863 -1656 11018
rect 35828 9167 35940 15204
rect 36058 9716 36158 15782
rect 36254 15507 36354 16103
rect 36249 15409 36255 15507
rect 36353 15409 36359 15507
rect 35828 9065 35833 9167
rect 35935 9065 35940 9167
rect 35828 9060 35940 9065
rect 36054 9395 36158 9716
rect 36254 9541 36354 15409
rect 36458 13717 36558 16322
rect 36451 13712 36561 13717
rect 36451 13612 36456 13712
rect 36556 13612 36561 13712
rect 36451 13607 36561 13612
rect 36249 9443 36255 9541
rect 36353 9443 36359 9541
rect 36254 9442 36354 9443
rect 36054 9390 36165 9395
rect 36054 9290 36060 9390
rect 36160 9290 36165 9390
rect 36054 9285 36165 9290
rect -1761 8765 -1755 8863
rect -1657 8765 -1651 8863
rect -11351 8460 -10749 8462
rect -8581 8460 -7979 8462
rect -7510 8460 -2607 8462
rect -12325 7873 -2607 8460
rect -12325 7871 -4183 7873
rect -12325 7860 -11351 7871
rect -10749 7862 -4183 7871
rect -10749 7860 -6351 7862
rect -11351 7263 -10749 7269
rect -8581 7851 -7979 7860
rect -8581 7243 -7979 7249
rect -6953 7853 -6351 7860
rect -6351 7251 -6332 7538
rect -3581 7862 -2607 7873
rect 35229 7738 35327 7743
rect -4183 7265 -3581 7271
rect 11362 7737 35328 7738
rect 11362 7639 35229 7737
rect 35327 7639 35328 7737
rect 11362 7638 35328 7639
rect -6953 7245 -6332 7251
rect -6932 7112 -6332 7245
rect 11362 7198 11462 7638
rect 35229 7633 35327 7638
rect 11362 7138 11382 7198
rect 11442 7138 11462 7198
rect -11324 7104 -10724 7110
rect -12309 6504 -11324 6560
rect -8544 7104 -7944 7110
rect -10724 6504 -8544 6560
rect -6956 7106 -6332 7112
rect -7720 6560 -6956 6562
rect -7944 6506 -6956 6560
rect -6356 6562 -6332 7106
rect -4176 7106 -3576 7112
rect -6356 6506 -4176 6562
rect 11362 7102 11462 7138
rect -3576 6506 -2591 6562
rect -7944 6504 -2591 6506
rect -12309 5962 -2591 6504
rect -12309 5960 -7650 5962
rect -12737 5567 -12731 5665
rect -12633 5567 -12627 5665
rect -12732 5566 -12632 5567
rect -12309 4926 -11709 5960
rect -12896 4326 -12890 4926
rect -12290 4326 -11709 4926
rect -12309 2848 -11709 4326
rect -9948 5696 -7198 5796
rect -9948 3640 -9848 5696
rect -7298 5478 -7198 5696
rect -3191 4928 -2591 5962
rect -2426 5665 -2322 5666
rect -2427 5567 -2421 5665
rect -2323 5567 -2317 5665
rect -2426 5228 -2322 5567
rect -2426 5226 8314 5228
rect -2426 5204 8366 5226
rect -2426 5144 8280 5204
rect 8340 5144 8366 5204
rect -2426 5126 8366 5144
rect -2426 5124 8314 5126
rect -3191 4328 -2610 4928
rect -2010 4328 -2004 4928
rect -10140 3637 -10040 3638
rect -10145 3539 -10139 3637
rect -10041 3539 -10035 3637
rect -9948 3540 -9374 3640
rect -9246 3638 -9146 3876
rect -8085 3644 -7987 3649
rect -7554 3644 -7454 3650
rect -8086 3643 -7554 3644
rect -10140 3350 -10040 3539
rect -10140 3238 -9986 3350
rect -9474 3254 -9374 3540
rect -9252 3538 -9246 3638
rect -9146 3538 -9140 3638
rect -8086 3545 -8085 3643
rect -7987 3545 -7554 3643
rect -8086 3544 -7554 3545
rect -5748 3640 -5648 3890
rect -5940 3637 -5840 3638
rect -8085 3539 -7987 3544
rect -7554 3538 -7454 3544
rect -5945 3539 -5939 3637
rect -5841 3539 -5835 3637
rect -5748 3540 -5174 3640
rect -5046 3638 -4946 3876
rect -3885 3644 -3787 3649
rect -3354 3644 -3254 3650
rect -3886 3643 -3354 3644
rect -7176 3254 -7174 3446
rect -5940 3238 -5840 3539
rect -5274 3446 -5174 3540
rect -5052 3538 -5046 3638
rect -4946 3538 -4940 3638
rect -3886 3545 -3885 3643
rect -3787 3545 -3354 3643
rect -3886 3544 -3354 3545
rect -3885 3539 -3787 3544
rect -3354 3538 -3254 3544
rect -5274 3254 -5176 3446
rect -12906 2248 -12900 2848
rect -12300 2248 -11709 2848
rect -13103 1529 -13097 1627
rect -12999 1529 -12993 1627
rect -13100 1528 -13000 1529
rect -12309 1222 -11709 2248
rect -10086 1474 -9986 3238
rect -3191 2850 -2591 4328
rect -3191 2250 -2600 2850
rect -2000 2250 -1994 2850
rect -7176 1474 -7076 1916
rect -10086 1374 -7076 1474
rect -6937 1224 -6335 1226
rect -4167 1224 -3565 1226
rect -3191 1224 -2591 2250
rect 36054 2238 36158 9285
rect 36458 6111 36558 13607
rect 36748 13581 36852 17048
rect 37297 16666 37897 18350
rect 39810 17674 39910 19730
rect 42460 19512 42560 19730
rect 46664 19432 46764 19730
rect 50792 18954 51393 19984
rect 50792 18354 51374 18954
rect 51974 18354 51980 18954
rect 39618 17671 39718 17672
rect 39613 17573 39619 17671
rect 39717 17573 39723 17671
rect 39810 17574 40384 17674
rect 40512 17672 40612 17910
rect 41673 17678 41771 17683
rect 42204 17678 42304 17684
rect 41672 17677 42204 17678
rect 39618 17384 39718 17573
rect 39618 17272 39772 17384
rect 40284 17288 40384 17574
rect 40506 17572 40512 17672
rect 40612 17572 40618 17672
rect 41672 17579 41673 17677
rect 41771 17579 42204 17677
rect 41672 17578 42204 17579
rect 44010 17674 44110 17924
rect 43818 17671 43918 17672
rect 41673 17573 41771 17578
rect 42204 17572 42304 17578
rect 43813 17573 43819 17671
rect 43917 17573 43923 17671
rect 44010 17574 44584 17674
rect 44712 17672 44812 17910
rect 45873 17678 45971 17683
rect 46404 17678 46504 17684
rect 45872 17677 46404 17678
rect 42582 17288 42584 17480
rect 43818 17272 43918 17573
rect 44484 17480 44584 17574
rect 44706 17572 44712 17672
rect 44812 17572 44818 17672
rect 45872 17579 45873 17677
rect 45971 17579 46404 17677
rect 45872 17578 46404 17579
rect 48210 17674 48310 17924
rect 48018 17671 48118 17672
rect 45873 17573 45971 17578
rect 46404 17572 46504 17578
rect 48013 17573 48019 17671
rect 48117 17573 48123 17671
rect 48210 17574 48784 17674
rect 48912 17672 49012 17910
rect 50073 17678 50171 17683
rect 50604 17678 50704 17684
rect 50072 17677 50604 17678
rect 44484 17288 44582 17480
rect 48018 17272 48118 17573
rect 48684 17288 48784 17574
rect 48906 17572 48912 17672
rect 49012 17572 49018 17672
rect 50072 17579 50073 17677
rect 50171 17579 50604 17677
rect 50072 17578 50604 17579
rect 50073 17573 50171 17578
rect 50604 17572 50704 17578
rect 36943 16380 36949 16666
rect 37235 16380 37897 16666
rect 37297 15248 37897 16380
rect 39672 15508 39772 17272
rect 50792 16876 51393 18354
rect 50792 16276 51384 16876
rect 51984 16276 51990 16876
rect 42582 15508 42682 15950
rect 46660 15508 46760 15844
rect 39292 15408 39298 15508
rect 39398 15408 46760 15508
rect 44725 15250 45327 15252
rect 47709 15250 48311 15252
rect 49817 15250 50419 15252
rect 50792 15250 51393 16276
rect 44268 15248 46396 15250
rect 46668 15248 51393 15250
rect 37297 14661 51393 15248
rect 37297 14648 49817 14661
rect 37297 14646 47259 14648
rect 37302 14478 47032 14646
rect 47709 14641 48311 14648
rect 37302 13942 47037 14478
rect 50419 14650 51393 14661
rect 52144 14738 52244 23614
rect 65088 18913 65188 18918
rect 65088 18823 65093 18913
rect 65183 18823 65188 18913
rect 65088 18818 65188 18823
rect 52380 15100 52480 15106
rect 64976 15100 65076 16422
rect 52480 15000 65076 15100
rect 52380 14994 52480 15000
rect 65083 14738 65193 14743
rect 50419 14648 51392 14650
rect 52144 14638 65088 14738
rect 65188 14638 65193 14738
rect 65083 14633 65193 14638
rect 49817 14053 50419 14059
rect 47709 14033 48311 14039
rect 37319 13832 47037 13942
rect 36743 13483 36749 13581
rect 36847 13483 36853 13581
rect 36748 13480 36852 13483
rect 37319 12842 37919 13832
rect 39248 13707 42430 13712
rect 39248 13617 39253 13707
rect 39343 13617 42430 13707
rect 39248 13612 42430 13617
rect 36732 12242 36738 12842
rect 37338 12242 37919 12842
rect 37319 10764 37919 12242
rect 39680 11556 39780 13612
rect 42330 13394 42430 13612
rect 46437 12844 47037 13832
rect 46437 12244 47018 12844
rect 47618 12244 47624 12844
rect 39488 11553 39588 11554
rect 39483 11455 39489 11553
rect 39587 11455 39593 11553
rect 39680 11456 40254 11556
rect 40382 11554 40482 11792
rect 41543 11560 41641 11565
rect 42074 11560 42174 11566
rect 41542 11559 42074 11560
rect 39488 11266 39588 11455
rect 39488 11154 39642 11266
rect 40154 11170 40254 11456
rect 40376 11454 40382 11554
rect 40482 11454 40488 11554
rect 41542 11461 41543 11559
rect 41641 11461 42074 11559
rect 41542 11460 42074 11461
rect 43880 11556 43980 11806
rect 43688 11553 43788 11554
rect 41543 11455 41641 11460
rect 42074 11454 42174 11460
rect 43683 11455 43689 11553
rect 43787 11455 43793 11553
rect 43880 11456 44454 11556
rect 44582 11554 44682 11792
rect 45743 11560 45841 11565
rect 46274 11560 46374 11566
rect 45742 11559 46274 11560
rect 42452 11170 42454 11362
rect 43688 11154 43788 11455
rect 44354 11362 44454 11456
rect 44576 11454 44582 11554
rect 44682 11454 44688 11554
rect 45742 11461 45743 11559
rect 45841 11461 46274 11559
rect 45742 11460 46274 11461
rect 45743 11455 45841 11460
rect 46274 11454 46374 11460
rect 44354 11170 44452 11362
rect 36722 10164 36728 10764
rect 37328 10164 37919 10764
rect 37319 9138 37919 10164
rect 39542 9390 39642 11154
rect 46437 10766 47037 12244
rect 46437 10166 47028 10766
rect 47628 10166 47634 10766
rect 42452 9390 42552 9832
rect 39004 9385 42552 9390
rect 39004 9295 39009 9385
rect 39099 9295 42552 9385
rect 39004 9290 42552 9295
rect 42691 9140 43293 9142
rect 45461 9140 46063 9142
rect 46437 9140 47037 10166
rect 38293 9138 38895 9140
rect 41063 9138 41665 9140
rect 42134 9138 47037 9140
rect 37319 8551 47037 9138
rect 37319 8549 45461 8551
rect 37319 8538 38293 8549
rect 38895 8540 45461 8549
rect 38895 8538 43293 8540
rect 38293 7941 38895 7947
rect 41063 8529 41665 8538
rect 41063 7921 41665 7927
rect 42691 8531 43293 8538
rect 46063 8540 47037 8551
rect 45461 7943 46063 7949
rect 42691 7923 43293 7929
rect 36990 7638 36996 7738
rect 37096 7638 47596 7738
rect 53050 7722 53150 7728
rect 38304 7420 38904 7426
rect 37319 6820 38304 6876
rect 41084 7420 41684 7426
rect 38904 6820 41084 6876
rect 42672 7422 43272 7428
rect 41908 6876 42672 6878
rect 41684 6822 42672 6876
rect 45452 7422 46052 7428
rect 43272 6822 45452 6878
rect 47496 7222 47596 7638
rect 49800 7700 53050 7722
rect 49800 7640 49822 7700
rect 49882 7640 53050 7700
rect 49800 7622 53050 7640
rect 53050 7616 53150 7622
rect 47494 7198 62432 7222
rect 47494 7138 62350 7198
rect 62410 7138 62432 7198
rect 47494 7122 62432 7138
rect 46052 6822 47037 6878
rect 41684 6820 47037 6822
rect 37319 6278 47037 6820
rect 37319 6276 41978 6278
rect 36453 6013 36459 6111
rect 36557 6013 36563 6111
rect 36458 6012 36558 6013
rect 37319 5242 37919 6276
rect 39048 6012 39054 6112
rect 39154 6107 46348 6112
rect 39154 6017 46253 6107
rect 46343 6017 46348 6107
rect 39154 6012 46348 6017
rect 36732 4642 36738 5242
rect 37338 4642 37919 5242
rect 37319 3164 37919 4642
rect 39680 3956 39780 6012
rect 42330 5794 42430 6012
rect 46437 5244 47037 6278
rect 48476 5981 48576 5982
rect 48471 5883 48477 5981
rect 48575 5883 48581 5981
rect 48476 5758 48576 5883
rect 48476 5736 49388 5758
rect 48476 5676 49306 5736
rect 49366 5676 49388 5736
rect 48476 5658 49388 5676
rect 53048 5604 53148 5610
rect 49924 5587 53048 5604
rect 49924 5527 49940 5587
rect 50000 5527 53048 5587
rect 49924 5504 53048 5527
rect 53048 5498 53148 5504
rect 46437 4644 47018 5244
rect 47618 4644 47624 5244
rect 52183 4956 52281 4961
rect 52183 4955 66110 4956
rect 52281 4936 66110 4955
rect 52281 4876 66026 4936
rect 66086 4876 66110 4936
rect 52281 4857 66110 4876
rect 52183 4856 66110 4857
rect 52183 4851 52281 4856
rect 39488 3953 39588 3954
rect 39483 3855 39489 3953
rect 39587 3855 39593 3953
rect 39680 3856 40254 3956
rect 40382 3954 40482 4192
rect 41543 3960 41641 3965
rect 42074 3960 42174 3966
rect 41542 3959 42074 3960
rect 39488 3666 39588 3855
rect 39488 3554 39642 3666
rect 40154 3570 40254 3856
rect 40376 3854 40382 3954
rect 40482 3854 40488 3954
rect 41542 3861 41543 3959
rect 41641 3861 42074 3959
rect 41542 3860 42074 3861
rect 43880 3956 43980 4206
rect 43688 3953 43788 3954
rect 41543 3855 41641 3860
rect 42074 3854 42174 3860
rect 43683 3855 43689 3953
rect 43787 3855 43793 3953
rect 43880 3856 44454 3956
rect 44582 3954 44682 4192
rect 45743 3960 45841 3965
rect 46274 3960 46374 3966
rect 45742 3959 46274 3960
rect 42452 3570 42454 3762
rect 43688 3554 43788 3855
rect 44354 3762 44454 3856
rect 44576 3854 44582 3954
rect 44682 3854 44688 3954
rect 45742 3861 45743 3959
rect 45841 3861 46274 3959
rect 45742 3860 46274 3861
rect 45743 3855 45841 3860
rect 46274 3854 46374 3860
rect 44354 3570 44452 3762
rect 36722 2564 36728 3164
rect 37328 2564 37919 3164
rect 36054 1789 36154 2238
rect 36049 1691 36055 1789
rect 36153 1691 36159 1789
rect 36054 1690 36154 1691
rect -2334 1625 -2234 1626
rect -2339 1527 -2333 1625
rect -2235 1527 -2229 1625
rect 37319 1538 37919 2564
rect 39542 1790 39642 3554
rect 46437 3166 47037 4644
rect 48482 3756 48582 3762
rect 48582 3736 49378 3756
rect 48582 3676 49302 3736
rect 49362 3676 49378 3736
rect 48582 3656 49378 3676
rect 48482 3650 48582 3656
rect 52181 3605 52283 3611
rect 50066 3587 52181 3604
rect 50066 3527 50082 3587
rect 50142 3527 52181 3587
rect 50066 3504 52181 3527
rect 52181 3497 52283 3503
rect 46437 2566 47028 3166
rect 47628 2566 47634 3166
rect 61918 2933 62248 2938
rect 61918 2843 62153 2933
rect 62243 2843 62248 2933
rect 53051 2834 53149 2839
rect 61918 2838 62248 2843
rect 61918 2834 62018 2838
rect 53051 2833 62018 2834
rect 53149 2735 62018 2833
rect 53051 2734 62018 2735
rect 53051 2729 53149 2734
rect 42452 1790 42552 2232
rect 39160 1690 39166 1790
rect 39266 1768 46374 1790
rect 39266 1708 46288 1768
rect 46348 1708 46374 1768
rect 39266 1690 46374 1708
rect 42691 1540 43293 1542
rect 45461 1540 46063 1542
rect 46437 1540 47037 2566
rect 52177 1672 52287 1678
rect 49806 1646 52177 1672
rect 49806 1586 49828 1646
rect 49888 1586 52177 1646
rect 49806 1562 52177 1586
rect 52177 1556 52287 1562
rect 38293 1538 38895 1540
rect 41063 1538 41665 1540
rect 42134 1538 47037 1540
rect -11335 1222 -10733 1224
rect -8565 1222 -7963 1224
rect -7494 1222 -2591 1224
rect -12309 635 -2591 1222
rect -12309 633 -4167 635
rect -12309 622 -11335 633
rect -10733 624 -4167 633
rect -10733 622 -6335 624
rect -11335 25 -10733 31
rect -8565 613 -7963 622
rect -8565 5 -7963 11
rect -6937 615 -6335 622
rect -3565 624 -2591 635
rect -2334 602 -2230 1527
rect 37319 951 47037 1538
rect 37319 949 45461 951
rect 37319 938 38293 949
rect -2334 582 8126 602
rect -2334 522 8042 582
rect 8102 522 8126 582
rect -2334 502 8126 522
rect -2334 500 -2234 502
rect 38895 940 45461 949
rect 38895 938 43293 940
rect 38293 341 38895 347
rect 41063 929 41665 938
rect 41063 321 41665 327
rect 42691 931 43293 938
rect 46063 940 47037 951
rect 45461 343 46063 349
rect 42691 323 43293 329
rect -4167 27 -3565 33
rect -6937 7 -6335 13
<< via3 >>
rect -1419 27642 -1349 27647
rect -1419 27583 -1414 27642
rect -1414 27583 -1354 27642
rect -1354 27583 -1349 27642
rect 47824 27564 48462 27680
rect 38288 26378 38888 27302
rect 41068 26378 41668 27302
rect 36734 24400 37334 25000
rect 36469 23607 36567 23705
rect 39509 23607 39607 23705
rect 42904 24440 43504 25040
rect 46576 24434 46676 24534
rect 36738 22324 37338 22924
rect 40402 23606 40502 23706
rect 41563 23613 41661 23711
rect 42094 23612 42194 23712
rect 42914 22312 43514 22912
rect 44725 20598 45327 21200
rect 49760 21600 49860 21700
rect 46405 21005 46503 21103
rect 47028 20532 47628 21132
rect 49808 20532 50408 21132
rect 52144 23614 52244 23714
rect 51794 20966 51894 21066
rect 36473 19731 36571 19829
rect 39078 19730 39178 19830
rect 36716 18350 37316 18950
rect -13471 10777 -13373 10875
rect -11340 13742 -10740 14342
rect -8560 13742 -7960 14342
rect -6972 13744 -6372 14344
rect -4192 13744 -3592 14344
rect -13107 12935 -13009 13033
rect -10574 12934 -10474 13034
rect -12906 11564 -12306 12164
rect -2396 12804 -2296 12904
rect -2626 11566 -2026 12166
rect -10155 10777 -10057 10875
rect -9262 10776 -9162 10876
rect -8101 10783 -8003 10881
rect -7570 10782 -7470 10882
rect -5955 10777 -5857 10875
rect -5062 10776 -4962 10876
rect -3901 10781 -3803 10879
rect -3370 10780 -3270 10880
rect -12916 9486 -12316 10086
rect -13099 8613 -13001 8711
rect -13303 3539 -13205 3637
rect -2616 9488 -2016 10088
rect -10504 8612 -10404 8712
rect 36255 15409 36353 15507
rect 36255 9443 36353 9541
rect -1755 8765 -1657 8863
rect -11351 7269 -10749 7871
rect -8581 7249 -7979 7851
rect -6953 7251 -6351 7853
rect -4183 7271 -3581 7873
rect 35229 7639 35327 7737
rect -11324 6504 -10724 7104
rect -8544 6504 -7944 7104
rect -6956 6506 -6356 7106
rect -4176 6506 -3576 7106
rect -12731 5567 -12633 5665
rect -12890 4326 -12290 4926
rect -2421 5567 -2323 5665
rect -2610 4328 -2010 4928
rect -10139 3539 -10041 3637
rect -9246 3538 -9146 3638
rect -8085 3545 -7987 3643
rect -7554 3544 -7454 3644
rect -5939 3539 -5841 3637
rect -5046 3538 -4946 3638
rect -3885 3545 -3787 3643
rect -3354 3544 -3254 3644
rect -12900 2248 -12300 2848
rect -13097 1529 -12999 1627
rect -2600 2250 -2000 2850
rect 51374 18354 51974 18954
rect 39619 17573 39717 17671
rect 40512 17572 40612 17672
rect 41673 17579 41771 17677
rect 42204 17578 42304 17678
rect 43819 17573 43917 17671
rect 44712 17572 44812 17672
rect 45873 17579 45971 17677
rect 46404 17578 46504 17678
rect 48019 17573 48117 17671
rect 48912 17572 49012 17672
rect 50073 17579 50171 17677
rect 50604 17578 50704 17678
rect 36949 16380 37235 16666
rect 51384 16276 51984 16876
rect 39298 15408 39398 15508
rect 47709 14039 48311 14641
rect 49817 14059 50419 14661
rect 52380 15000 52480 15100
rect 36749 13483 36847 13581
rect 36738 12242 37338 12842
rect 47018 12244 47618 12844
rect 39489 11455 39587 11553
rect 40382 11454 40482 11554
rect 41543 11461 41641 11559
rect 42074 11460 42174 11560
rect 43689 11455 43787 11553
rect 44582 11454 44682 11554
rect 45743 11461 45841 11559
rect 46274 11460 46374 11560
rect 36728 10164 37328 10764
rect 47028 10166 47628 10766
rect 38293 7947 38895 8549
rect 41063 7927 41665 8529
rect 42691 7929 43293 8531
rect 45461 7949 46063 8551
rect 36996 7638 37096 7738
rect 38304 6820 38904 7420
rect 41084 6820 41684 7420
rect 42672 6822 43272 7422
rect 45452 6822 46052 7422
rect 53050 7622 53150 7722
rect 36459 6013 36557 6111
rect 39054 6012 39154 6112
rect 36738 4642 37338 5242
rect 48477 5883 48575 5981
rect 53048 5504 53148 5604
rect 47018 4644 47618 5244
rect 52183 4857 52281 4955
rect 39489 3855 39587 3953
rect 40382 3854 40482 3954
rect 41543 3861 41641 3959
rect 42074 3860 42174 3960
rect 43689 3855 43787 3953
rect 44582 3854 44682 3954
rect 45743 3861 45841 3959
rect 46274 3860 46374 3960
rect 36728 2564 37328 3164
rect 36055 1691 36153 1789
rect -2333 1527 -2235 1625
rect 48482 3656 48582 3756
rect 52181 3503 52283 3605
rect 47028 2566 47628 3166
rect 53051 2735 53149 2833
rect 39166 1690 39266 1790
rect 52177 1562 52287 1672
rect -11335 31 -10733 633
rect -8565 11 -7963 613
rect -6937 13 -6335 615
rect -4167 33 -3565 635
rect 38293 347 38895 949
rect 41063 327 41665 929
rect 42691 329 43293 931
rect 45461 349 46063 951
<< metal4 >>
rect 33530 27680 55572 28340
rect -1420 27647 -1348 27648
rect -1420 27583 -1419 27647
rect -1349 27583 -1348 27647
rect -1420 27582 -1348 27583
rect 33530 27564 47824 27680
rect 48462 27564 55572 27680
rect 33530 27540 55572 27564
rect 38287 27302 38889 27303
rect 38287 26378 38288 27302
rect 38888 26378 38889 27302
rect 38287 26377 38889 26378
rect 41067 27302 41669 27303
rect 41067 26378 41068 27302
rect 41668 26378 41669 27302
rect 41067 26377 41669 26378
rect 38288 25826 38888 26377
rect 41068 25816 41668 26377
rect 39530 25634 46676 25734
rect 39530 25280 39630 25634
rect 36733 25000 37335 25001
rect 36733 24400 36734 25000
rect 37334 24400 37896 25000
rect 41418 24614 41958 24714
rect 36733 24399 37335 24400
rect 41562 23711 41662 23712
rect 40401 23706 40503 23707
rect 36468 23705 40402 23706
rect 36468 23607 36469 23705
rect 36567 23607 39509 23705
rect 39607 23607 40402 23705
rect 36468 23606 40402 23607
rect 40502 23606 40503 23706
rect 40401 23605 40503 23606
rect 41562 23613 41563 23711
rect 41661 23613 41662 23711
rect 41562 23212 41662 23613
rect 36737 22924 37339 22925
rect 36737 22324 36738 22924
rect 37338 22324 37888 22924
rect 36737 22323 37339 22324
rect 39512 21694 39612 22074
rect 41858 21694 41958 24614
rect 42094 23714 42194 25634
rect 42903 25040 43505 25041
rect 42312 24440 42904 25040
rect 43504 24440 43505 25040
rect 46576 24535 46676 25634
rect 42903 24439 43505 24440
rect 46575 24534 46677 24535
rect 46575 24434 46576 24534
rect 46676 24434 46677 24534
rect 46575 24433 46677 24434
rect 52143 23714 52245 23715
rect 42094 23713 52144 23714
rect 42093 23712 52144 23713
rect 42093 23612 42094 23712
rect 42194 23614 52144 23712
rect 52244 23614 52245 23714
rect 42194 23612 42195 23614
rect 52143 23613 52245 23614
rect 42093 23611 42195 23612
rect 42913 22912 43515 22913
rect 42302 22312 42914 22912
rect 43514 22312 43515 22912
rect 42913 22311 43515 22312
rect 49759 21700 49861 21701
rect 49759 21694 49760 21700
rect 39512 21600 49760 21694
rect 49860 21694 49861 21700
rect 52380 21694 52480 21696
rect 49860 21600 52480 21694
rect 39512 21594 52480 21600
rect 38292 20888 42556 21370
rect 38292 20576 38496 20888
rect 42366 20598 42556 20888
rect 44724 21200 45328 21201
rect 44724 20598 44725 21200
rect 45327 20598 45328 21200
rect 47027 21132 47629 21133
rect 42366 20597 45328 20598
rect 46404 21103 46504 21104
rect 46404 21005 46405 21103
rect 46503 21005 46504 21103
rect 42366 20576 45327 20597
rect 38292 20026 45327 20576
rect 39077 19830 39179 19831
rect 36472 19829 39078 19830
rect 36472 19731 36473 19829
rect 36571 19731 39078 19829
rect 36472 19730 39078 19731
rect 39178 19730 39179 19830
rect 39077 19729 39179 19730
rect 46404 19700 46504 21005
rect 47027 20532 47028 21132
rect 47628 20532 47629 21132
rect 47027 20531 47629 20532
rect 49807 21132 50409 21133
rect 49807 20532 49808 21132
rect 50408 20532 50409 21132
rect 51793 21066 51895 21067
rect 51793 20966 51794 21066
rect 51894 20966 52248 21066
rect 51793 20965 51895 20966
rect 49807 20531 50409 20532
rect 47028 19970 47628 20531
rect 49808 19980 50408 20531
rect 39640 19600 50704 19700
rect 39640 19246 39740 19600
rect 36715 18950 37317 18951
rect 36715 18350 36716 18950
rect 37316 18350 37888 18950
rect 41528 18580 42068 18680
rect 36715 18349 37317 18350
rect 41672 17677 41772 17678
rect 40511 17672 40613 17673
rect 39618 17671 40512 17672
rect 39618 17573 39619 17671
rect 39717 17573 40512 17671
rect 39618 17572 40512 17573
rect 40612 17572 40613 17672
rect 40511 17571 40613 17572
rect 41672 17579 41673 17677
rect 41771 17579 41772 17677
rect 41672 17178 41772 17579
rect 36948 16666 37236 16667
rect 36948 16380 36949 16666
rect 37235 16380 37753 16666
rect 36948 16379 37236 16380
rect 39622 15660 39722 16040
rect 41968 15660 42068 18580
rect 42204 17679 42304 19600
rect 43840 19246 43940 19600
rect 45728 18580 46268 18680
rect 42203 17678 42305 17679
rect 42203 17578 42204 17678
rect 42304 17578 42305 17678
rect 45872 17677 45972 17678
rect 44711 17672 44813 17673
rect 42203 17577 42305 17578
rect 43818 17671 44712 17672
rect 43818 17573 43819 17671
rect 43917 17573 44712 17671
rect 43818 17572 44712 17573
rect 44812 17572 44813 17672
rect 44711 17571 44813 17572
rect 45872 17579 45873 17677
rect 45971 17579 45972 17677
rect 45872 17178 45972 17579
rect 43822 15660 43922 16040
rect 46168 15660 46268 18580
rect 46404 17679 46504 19600
rect 48040 19246 48140 19600
rect 49928 18580 50468 18680
rect 46403 17678 46505 17679
rect 46403 17578 46404 17678
rect 46504 17578 46505 17678
rect 50072 17677 50172 17678
rect 48911 17672 49013 17673
rect 46403 17577 46505 17578
rect 48018 17671 48912 17672
rect 48018 17573 48019 17671
rect 48117 17573 48912 17671
rect 48018 17572 48912 17573
rect 49012 17572 49013 17672
rect 48911 17571 49013 17572
rect 50072 17579 50073 17677
rect 50171 17579 50172 17677
rect 50072 17178 50172 17579
rect 48022 15660 48122 16040
rect 50368 15660 50468 18580
rect 50604 17679 50704 19600
rect 51373 18954 51975 18955
rect 50802 18354 51374 18954
rect 51974 18354 51975 18954
rect 51373 18353 51975 18354
rect 50603 17678 50705 17679
rect 50603 17578 50604 17678
rect 50704 17578 50705 17678
rect 50603 17577 50705 17578
rect 51383 16876 51985 16877
rect 50812 16276 51384 16876
rect 51984 16276 51985 16876
rect 51383 16275 51985 16276
rect 52148 15660 52248 20966
rect 39622 15560 52248 15660
rect 39297 15508 39399 15509
rect 36254 15507 39298 15508
rect 36254 15409 36255 15507
rect 36353 15409 39298 15507
rect 36254 15408 39298 15409
rect 39398 15408 39399 15508
rect 39297 15407 39399 15408
rect 47610 15111 48410 15242
rect 37509 14804 48410 15111
rect 37509 14348 37816 14804
rect 45494 14768 46046 14804
rect 47610 14641 48410 14804
rect 47610 14348 47709 14641
rect -6973 14344 -6371 14345
rect -11341 14342 -10739 14343
rect -11341 13742 -11340 14342
rect -10740 13742 -10739 14342
rect -11341 13741 -10739 13742
rect -8561 14342 -7959 14343
rect -8561 13742 -8560 14342
rect -7960 13742 -7959 14342
rect -6973 13744 -6972 14344
rect -6372 13744 -6371 14344
rect -6973 13743 -6371 13744
rect -4193 14344 -3591 14345
rect -4193 13744 -4192 14344
rect -3592 13744 -3591 14344
rect 37509 14041 47709 14348
rect -4193 13743 -3591 13744
rect 47610 14039 47709 14041
rect 48311 14039 48410 14641
rect -8561 13741 -7959 13742
rect -11340 13190 -10740 13741
rect -8560 13180 -7960 13741
rect -6972 13182 -6372 13743
rect -4192 13192 -3592 13743
rect 47610 13732 48410 14039
rect 49718 14661 50518 15252
rect 52380 15101 52480 21594
rect 52379 15100 52481 15101
rect 52379 15000 52380 15100
rect 52480 15000 52481 15100
rect 52379 14999 52481 15000
rect 49718 14059 49817 14661
rect 50419 14059 50518 14661
rect 49718 13732 50518 14059
rect 36748 13581 46374 13582
rect 36748 13483 36749 13581
rect 36847 13483 46374 13581
rect 36748 13482 46374 13483
rect 39510 13128 39610 13482
rect -10575 13034 -10473 13035
rect -13108 13033 -10574 13034
rect -13108 12935 -13107 13033
rect -13009 12935 -10574 13033
rect -13108 12934 -10574 12935
rect -10474 12934 -10473 13034
rect -10575 12933 -10473 12934
rect -2397 12904 -2295 12905
rect -10134 12804 -2396 12904
rect -2296 12804 -2295 12904
rect -10134 12450 -10034 12804
rect -12907 12164 -12305 12165
rect -12907 11564 -12906 12164
rect -12306 11564 -11734 12164
rect -8246 11784 -7706 11884
rect -12907 11563 -12305 11564
rect -8102 10881 -8002 10882
rect -9263 10876 -9161 10877
rect -13472 10875 -9262 10876
rect -13472 10777 -13471 10875
rect -13373 10777 -10155 10875
rect -10057 10777 -9262 10875
rect -13472 10776 -9262 10777
rect -9162 10776 -9161 10876
rect -9263 10775 -9161 10776
rect -8102 10783 -8101 10881
rect -8003 10783 -8002 10881
rect -8102 10382 -8002 10783
rect -12917 10086 -12315 10087
rect -12917 9486 -12916 10086
rect -12316 9486 -11744 10086
rect -12917 9485 -12315 9486
rect -10152 8864 -10052 9244
rect -7806 8864 -7706 11784
rect -7570 10883 -7470 12804
rect -5934 12450 -5834 12804
rect -4046 11784 -3506 11884
rect -7571 10882 -7469 10883
rect -7571 10782 -7570 10882
rect -7470 10782 -7469 10882
rect -3902 10879 -3802 10880
rect -5063 10876 -4961 10877
rect -7571 10781 -7469 10782
rect -5956 10875 -5062 10876
rect -5956 10777 -5955 10875
rect -5857 10777 -5062 10875
rect -5956 10776 -5062 10777
rect -4962 10776 -4961 10876
rect -5063 10775 -4961 10776
rect -3902 10781 -3901 10879
rect -3803 10781 -3802 10879
rect -3902 10382 -3802 10781
rect -5952 8864 -5852 9244
rect -3606 8864 -3506 11784
rect -3370 10881 -3270 12804
rect -2397 12803 -2295 12804
rect 36737 12842 37339 12843
rect 36737 12242 36738 12842
rect 37338 12242 37910 12842
rect 41398 12462 41938 12562
rect 36737 12241 37339 12242
rect -2627 12166 -2025 12167
rect -3198 11566 -2626 12166
rect -2026 11566 -2025 12166
rect -2627 11565 -2025 11566
rect 41542 11559 41642 11560
rect 40381 11554 40483 11555
rect 39488 11553 40382 11554
rect 39488 11455 39489 11553
rect 39587 11455 40382 11553
rect 39488 11454 40382 11455
rect 40482 11454 40483 11554
rect 40381 11453 40483 11454
rect 41542 11461 41543 11559
rect 41641 11461 41642 11559
rect 41542 11060 41642 11461
rect -3371 10880 -3269 10881
rect -3371 10780 -3370 10880
rect -3270 10780 -3269 10880
rect -3371 10779 -3269 10780
rect 36727 10764 37329 10765
rect 36727 10164 36728 10764
rect 37328 10164 37900 10764
rect 36727 10163 37329 10164
rect -2617 10088 -2015 10089
rect -3188 9488 -2616 10088
rect -2016 9488 -2015 10088
rect 39492 9542 39592 9922
rect 41838 9542 41938 12462
rect 42074 11561 42174 13482
rect 43710 13128 43810 13482
rect 45598 12462 46138 12562
rect 42073 11560 42175 11561
rect 42073 11460 42074 11560
rect 42174 11460 42175 11560
rect 45742 11559 45842 11560
rect 44581 11554 44683 11555
rect 42073 11459 42175 11460
rect 43688 11553 44582 11554
rect 43688 11455 43689 11553
rect 43787 11455 44582 11553
rect 43688 11454 44582 11455
rect 44682 11454 44683 11554
rect 44581 11453 44683 11454
rect 45742 11461 45743 11559
rect 45841 11461 45842 11559
rect 45742 11060 45842 11461
rect 43692 9542 43792 9922
rect 46038 9542 46138 12462
rect 46274 11561 46374 13482
rect 47017 12844 47619 12845
rect 46446 12244 47018 12844
rect 47618 12244 47619 12844
rect 47017 12243 47619 12244
rect 46273 11560 46375 11561
rect 46273 11460 46274 11560
rect 46374 11556 46375 11560
rect 46374 11460 53150 11556
rect 46273 11459 53150 11460
rect 46274 11456 53150 11459
rect 47027 10766 47629 10767
rect 46456 10166 47028 10766
rect 47628 10166 47629 10766
rect 47027 10165 47629 10166
rect -2617 9487 -2015 9488
rect 36254 9541 52282 9542
rect 36254 9443 36255 9541
rect 36353 9443 52282 9541
rect 36254 9442 52282 9443
rect -10152 8863 -1656 8864
rect -10152 8765 -1755 8863
rect -1657 8765 -1656 8863
rect -10152 8764 -1656 8765
rect -10505 8712 -10403 8713
rect -13100 8711 -10504 8712
rect -13100 8613 -13099 8711
rect -13001 8613 -10504 8711
rect -13100 8612 -10504 8613
rect -10404 8612 -10403 8712
rect -10505 8611 -10403 8612
rect 38293 8550 38895 9131
rect 38292 8549 38896 8550
rect -11351 7872 -10749 8453
rect -11352 7871 -10748 7872
rect -11352 7269 -11351 7871
rect -10749 7269 -10748 7871
rect -8581 7852 -7979 8423
rect -6953 7854 -6351 8425
rect -4183 7874 -3581 8455
rect 38292 7947 38293 8549
rect 38895 7947 38896 8549
rect 41063 8530 41665 9101
rect 42691 8532 43293 9103
rect 45461 8552 46063 9133
rect 45460 8551 46064 8552
rect 42690 8531 43294 8532
rect 38292 7946 38896 7947
rect 41062 8529 41666 8530
rect -4184 7873 -3580 7874
rect -6954 7853 -6350 7854
rect -11352 7268 -10748 7269
rect -8582 7851 -7978 7852
rect -11306 7105 -10754 7268
rect -8582 7249 -8581 7851
rect -7979 7519 -7978 7851
rect -7979 7249 -7955 7519
rect -6954 7517 -6953 7853
rect -8582 7248 -7955 7249
rect -8517 7105 -7955 7248
rect -6956 7251 -6953 7517
rect -6351 7251 -6350 7853
rect -4184 7271 -4183 7873
rect -3581 7498 -3580 7873
rect 36995 7738 37097 7739
rect 35228 7737 36996 7738
rect 35228 7639 35229 7737
rect 35327 7639 36996 7737
rect 35228 7638 36996 7639
rect 37096 7638 37097 7738
rect 36995 7637 37097 7638
rect -3581 7271 -3576 7498
rect 38304 7421 38856 7946
rect 41062 7927 41063 8529
rect 41665 7927 41666 8529
rect 42690 7929 42691 8531
rect 43293 7929 43294 8531
rect 45460 7949 45461 8551
rect 46063 7949 46064 8551
rect 45460 7948 46064 7949
rect 42690 7928 43294 7929
rect 41062 7926 41666 7927
rect 41084 7421 41646 7926
rect 42710 7423 43272 7928
rect 45500 7423 46052 7948
rect 42671 7422 43273 7423
rect -4184 7270 -3576 7271
rect -6956 7250 -6350 7251
rect -6956 7107 -6394 7250
rect -4128 7107 -3576 7270
rect 38303 7420 38905 7421
rect -6957 7106 -6355 7107
rect -11325 7104 -10723 7105
rect -11325 6504 -11324 7104
rect -10724 6504 -10723 7104
rect -11325 6503 -10723 6504
rect -8545 7104 -7943 7105
rect -8545 6504 -8544 7104
rect -7944 6504 -7943 7104
rect -6957 6506 -6956 7106
rect -6356 6506 -6355 7106
rect -6957 6505 -6355 6506
rect -4177 7106 -3575 7107
rect -4177 6506 -4176 7106
rect -3576 6506 -3575 7106
rect 38303 6820 38304 7420
rect 38904 6820 38905 7420
rect 38303 6819 38905 6820
rect 41083 7420 41685 7421
rect 41083 6820 41084 7420
rect 41684 6820 41685 7420
rect 42671 6822 42672 7422
rect 43272 6822 43273 7422
rect 42671 6821 43273 6822
rect 45451 7422 46053 7423
rect 45451 6822 45452 7422
rect 46052 6822 46053 7422
rect 45451 6821 46053 6822
rect 41083 6819 41685 6820
rect -4177 6505 -3575 6506
rect -8545 6503 -7943 6504
rect -11324 5952 -10724 6503
rect -8544 5942 -7944 6503
rect -6956 5944 -6356 6505
rect -4176 5954 -3576 6505
rect 38304 6268 38904 6819
rect 41084 6258 41684 6819
rect 42672 6260 43272 6821
rect 45452 6270 46052 6821
rect 39053 6112 39155 6113
rect 36458 6111 39054 6112
rect 36458 6013 36459 6111
rect 36557 6013 39054 6111
rect 36458 6012 39054 6013
rect 39154 6012 39155 6112
rect 39053 6011 39155 6012
rect 39510 5981 48576 5982
rect 39510 5883 48477 5981
rect 48575 5883 48576 5981
rect 39510 5882 48576 5883
rect -12732 5665 -2322 5666
rect -12732 5567 -12731 5665
rect -12633 5567 -2421 5665
rect -2323 5567 -2322 5665
rect -12732 5566 -2322 5567
rect -10118 5212 -10018 5566
rect -12891 4926 -12289 4927
rect -12891 4326 -12890 4926
rect -12290 4326 -11718 4926
rect -8230 4546 -7690 4646
rect -12891 4325 -12289 4326
rect -8086 3643 -7986 3644
rect -9247 3638 -9145 3639
rect -13304 3637 -9246 3638
rect -13304 3539 -13303 3637
rect -13205 3539 -10139 3637
rect -10041 3539 -9246 3637
rect -13304 3538 -9246 3539
rect -9146 3538 -9145 3638
rect -9247 3537 -9145 3538
rect -8086 3545 -8085 3643
rect -7987 3545 -7986 3643
rect -8086 3144 -7986 3545
rect -12901 2848 -12299 2849
rect -12901 2248 -12900 2848
rect -12300 2248 -11728 2848
rect -12901 2247 -12299 2248
rect -10136 1628 -10036 2006
rect -13098 1627 -9512 1628
rect -13098 1529 -13097 1627
rect -12999 1626 -9512 1627
rect -7790 1626 -7690 4546
rect -7554 3645 -7454 5566
rect -5918 5212 -5818 5566
rect -4030 4546 -3490 4646
rect -7555 3644 -7453 3645
rect -7555 3544 -7554 3644
rect -7454 3544 -7453 3644
rect -3886 3643 -3786 3644
rect -5047 3638 -4945 3639
rect -7555 3543 -7453 3544
rect -5940 3637 -5046 3638
rect -5940 3539 -5939 3637
rect -5841 3539 -5046 3637
rect -5940 3538 -5046 3539
rect -4946 3538 -4945 3638
rect -5047 3537 -4945 3538
rect -3886 3545 -3885 3643
rect -3787 3545 -3786 3643
rect -3886 3144 -3786 3545
rect -5936 1626 -5836 2006
rect -3590 1626 -3490 4546
rect -3354 3645 -3254 5566
rect 39510 5528 39610 5882
rect 36737 5242 37339 5243
rect -2611 4928 -2009 4929
rect -3182 4328 -2610 4928
rect -2010 4328 -2009 4928
rect 36737 4642 36738 5242
rect 37338 4642 37910 5242
rect 41398 4862 41938 4962
rect 36737 4641 37339 4642
rect -2611 4327 -2009 4328
rect 41542 3959 41642 3960
rect 40381 3954 40483 3955
rect 39488 3953 40382 3954
rect 39488 3855 39489 3953
rect 39587 3855 40382 3953
rect 39488 3854 40382 3855
rect 40482 3854 40483 3954
rect 40381 3853 40483 3854
rect 41542 3861 41543 3959
rect 41641 3861 41642 3959
rect -3355 3644 -3253 3645
rect -3355 3544 -3354 3644
rect -3254 3544 -3253 3644
rect -3355 3543 -3253 3544
rect 41542 3460 41642 3861
rect 36727 3164 37329 3165
rect -2601 2850 -1999 2851
rect -3172 2250 -2600 2850
rect -2000 2250 -1999 2850
rect 36727 2564 36728 3164
rect 37328 2564 37900 3164
rect 36727 2563 37329 2564
rect -2601 2249 -1999 2250
rect 39492 1942 39592 2322
rect 41838 1942 41938 4862
rect 42074 3961 42174 5882
rect 43710 5528 43810 5882
rect 45598 4862 46138 4962
rect 42073 3960 42175 3961
rect 42073 3860 42074 3960
rect 42174 3860 42175 3960
rect 45742 3959 45842 3960
rect 44581 3954 44683 3955
rect 42073 3859 42175 3860
rect 43688 3953 44582 3954
rect 43688 3855 43689 3953
rect 43787 3855 44582 3953
rect 43688 3854 44582 3855
rect 44682 3854 44683 3954
rect 44581 3853 44683 3854
rect 45742 3861 45743 3959
rect 45841 3861 45842 3959
rect 45742 3460 45842 3861
rect 43692 1942 43792 2322
rect 46038 1942 46138 4862
rect 46274 3961 46374 5882
rect 47017 5244 47619 5245
rect 46446 4644 47018 5244
rect 47618 4644 47619 5244
rect 47017 4643 47619 4644
rect 52182 4955 52282 9442
rect 53050 7723 53150 11456
rect 53049 7722 53151 7723
rect 53049 7622 53050 7722
rect 53150 7622 53151 7722
rect 53049 7621 53151 7622
rect 53050 5605 53150 7621
rect 53047 5604 53150 5605
rect 53047 5504 53048 5604
rect 53148 5504 53150 5604
rect 53047 5503 53150 5504
rect 52182 4857 52183 4955
rect 52281 4857 52282 4955
rect 52182 4087 52282 4857
rect 46273 3960 46375 3961
rect 46273 3860 46274 3960
rect 46374 3860 46375 3960
rect 46273 3859 46375 3860
rect 48481 3756 48583 3757
rect 48481 3656 48482 3756
rect 48582 3656 48583 3756
rect 48481 3655 48583 3656
rect 47027 3166 47629 3167
rect 46456 2566 47028 3166
rect 47628 2566 47629 3166
rect 47027 2565 47629 2566
rect 48482 1942 48582 3655
rect 52181 3606 52283 4087
rect 52180 3605 52284 3606
rect 52180 3503 52181 3605
rect 52283 3503 52284 3605
rect 52180 3502 52284 3503
rect 39492 1842 48582 1942
rect 52181 1897 52283 3502
rect 53050 2833 53150 5503
rect 53050 2735 53051 2833
rect 53149 2735 53150 2833
rect 53050 2734 53150 2735
rect 39165 1790 39267 1791
rect 36054 1789 39166 1790
rect 36054 1691 36055 1789
rect 36153 1691 39166 1789
rect 36054 1690 39166 1691
rect 39266 1690 39267 1790
rect 39165 1689 39267 1690
rect 52177 1673 52287 1897
rect 52176 1672 52288 1673
rect -12999 1625 -2234 1626
rect -12999 1529 -2333 1625
rect -13098 1528 -2333 1529
rect -10136 1527 -2333 1528
rect -2235 1527 -2234 1625
rect 52176 1562 52177 1672
rect 52287 1562 52288 1672
rect 52176 1561 52288 1562
rect -10136 1526 -2234 1527
rect -11350 633 -10550 1226
rect -11350 31 -11335 633
rect -10733 140 -10550 633
rect -8608 613 -7937 1231
rect -8608 140 -8565 613
rect -10733 31 -8565 140
rect -11350 11 -8565 31
rect -7963 140 -7937 613
rect -6990 615 -6317 1232
rect -6990 140 -6937 615
rect -7963 13 -6937 140
rect -6335 140 -6317 615
rect -4211 635 -3518 1252
rect -4211 140 -4167 635
rect -6335 33 -4167 140
rect -3565 140 -3518 635
rect 38202 949 39002 1544
rect 38202 347 38293 949
rect 38895 347 39002 949
rect 38202 140 39002 347
rect 40960 929 41760 1544
rect 40960 327 41063 929
rect 41665 327 41760 929
rect 40960 140 41760 327
rect 42596 931 43396 1544
rect 42596 329 42691 931
rect 43293 329 43396 931
rect 42596 140 43396 329
rect 45364 951 46164 1552
rect 45364 349 45461 951
rect 46063 349 46164 951
rect 45364 140 46164 349
rect -3565 33 378 140
rect -6335 13 378 33
rect -7963 11 378 13
rect -11350 -660 378 11
rect 34882 -660 90192 140
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_to_se_converter
timestamp 1624127230
transform 1 0 -8594 0 1 924
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_6 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_to_se_converter
timestamp 1624127230
transform 1 0 -10632 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_7
timestamp 1624127230
transform 1 0 -8632 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_4 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_to_se_converter
timestamp 1624127230
transform -1 0 -11077 0 1 924
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_4 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_to_se_converter
timestamp 1624127230
transform 1 0 -11958 0 1 2542
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_3
timestamp 1624127230
transform -1 0 -6306 0 1 926
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_9
timestamp 1624127230
transform 1 0 -6432 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_8
timestamp 1624127230
transform 1 0 -4432 0 1 2546
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_7
timestamp 1624127230
transform 1 0 -3823 0 1 926
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_7
timestamp 1624127230
transform -1 0 -2942 0 1 2544
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_5
timestamp 1624127230
transform 1 0 -10632 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_5
timestamp 1624127230
transform 1 0 -11958 0 1 4646
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_4
timestamp 1624127230
transform 1 0 -8632 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_5
timestamp 1624127230
transform -1 0 -11077 0 1 6260
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_1
timestamp 1624127230
transform 1 0 -8594 0 1 6260
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_10
timestamp 1624127230
transform 1 0 -6432 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_2
timestamp 1624127230
transform -1 0 -6306 0 1 6262
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_11
timestamp 1624127230
transform 1 0 -4432 0 1 4646
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_6
timestamp 1624127230
transform 1 0 -3823 0 1 6262
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_6
timestamp 1624127230
transform -1 0 -2942 0 1 4648
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_23
timestamp 1624127230
transform -1 0 -11093 0 1 8162
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_22
timestamp 1624127230
transform 1 0 -11974 0 1 9780
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_46
timestamp 1624127230
transform 1 0 -10648 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_22
timestamp 1624127230
transform 1 0 -8610 0 1 8162
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_42
timestamp 1624127230
transform 1 0 -8648 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_23
timestamp 1624127230
transform -1 0 -6322 0 1 8164
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_43
timestamp 1624127230
transform 1 0 -6448 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_22
timestamp 1624127230
transform 1 0 -3839 0 1 8164
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_40
timestamp 1624127230
transform 1 0 -4448 0 1 9784
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_20
timestamp 1624127230
transform -1 0 -2958 0 1 9782
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_23
timestamp 1624127230
transform 1 0 -11974 0 1 11884
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_47
timestamp 1624127230
transform 1 0 -10648 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_44
timestamp 1624127230
transform 1 0 -8648 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_21
timestamp 1624127230
transform -1 0 -11093 0 1 13498
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_20
timestamp 1624127230
transform 1 0 -8610 0 1 13498
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_45
timestamp 1624127230
transform 1 0 -6448 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_21
timestamp 1624127230
transform -1 0 -6322 0 1 13500
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_41
timestamp 1624127230
transform 1 0 -4448 0 1 11884
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_20
timestamp 1624127230
transform 1 0 -3839 0 1 13500
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_21
timestamp 1624127230
transform -1 0 -2958 0 1 11886
box -350 -900 244 900
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624127230
transform -1 0 -7834 0 1 15218
box -38 -48 314 592
use txgate  txgate_5 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/txgate
timestamp 1624127230
transform 1 0 -84715 0 1 -42708
box 74185 57360 76542 59116
use txgate  txgate_4
timestamp 1624127230
transform 1 0 -87315 0 1 -42708
box 74185 57360 76542 59116
use diff_fold_casc_ota  diff_fold_casc_ota_0 ~/ee272b/ee272b_mixed_signal_mmwave_accelerator/layouts/diff_fold_casc_ota
timestamp 1624135731
transform 1 0 10950 0 1 26540
box -12400 -27258 25000 1800
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_19
timestamp 1624127230
transform -1 0 38551 0 1 1240
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_38
timestamp 1624127230
transform 1 0 38996 0 1 2862
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_18
timestamp 1624127230
transform 1 0 37670 0 1 2858
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_35
timestamp 1624127230
transform 1 0 40996 0 1 2862
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_19
timestamp 1624127230
transform 1 0 41034 0 1 1240
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_18
timestamp 1624127230
transform -1 0 43322 0 1 1242
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_34
timestamp 1624127230
transform 1 0 43196 0 1 2862
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_18
timestamp 1624127230
transform 1 0 45805 0 1 1242
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_32
timestamp 1624127230
transform 1 0 45196 0 1 2862
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_16
timestamp 1624127230
transform -1 0 46686 0 1 2860
box -350 -900 244 900
use txgate  txgate_6
timestamp 1624127230
transform 1 0 -25531 0 1 -56596
box 74185 57360 76542 59116
use txgate  txgate_1
timestamp 1624127230
transform 1 0 -25531 0 1 -54506
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_19
timestamp 1624127230
transform 1 0 37670 0 1 4962
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_39
timestamp 1624127230
transform 1 0 38996 0 1 4962
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_17
timestamp 1624127230
transform -1 0 38551 0 1 6576
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_36
timestamp 1624127230
transform 1 0 40996 0 1 4962
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_16
timestamp 1624127230
transform 1 0 41034 0 1 6576
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_37
timestamp 1624127230
transform 1 0 43196 0 1 4962
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_17
timestamp 1624127230
transform -1 0 43322 0 1 6578
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_33
timestamp 1624127230
transform 1 0 45196 0 1 4962
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_16
timestamp 1624127230
transform 1 0 45805 0 1 6578
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_17
timestamp 1624127230
transform -1 0 46686 0 1 4964
box -350 -900 244 900
use txgate  txgate_0
timestamp 1624127230
transform 1 0 -25531 0 1 -52506
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_12
timestamp 1624127230
transform -1 0 38551 0 1 8840
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_25
timestamp 1624127230
transform 1 0 38996 0 1 10462
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_12
timestamp 1624127230
transform 1 0 37670 0 1 10458
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_12
timestamp 1624127230
transform 1 0 41034 0 1 8840
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_27
timestamp 1624127230
transform 1 0 40996 0 1 10462
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_13
timestamp 1624127230
transform -1 0 43322 0 1 8842
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_28
timestamp 1624127230
transform 1 0 43196 0 1 10462
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_13
timestamp 1624127230
transform 1 0 45805 0 1 8842
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_30
timestamp 1624127230
transform 1 0 45196 0 1 10462
box -950 -900 838 900
use txgate  txgate_7
timestamp 1624127230
transform 1 0 -25531 0 1 -50542
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_15
timestamp 1624127230
transform -1 0 46686 0 1 10460
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_24
timestamp 1624127230
transform 1 0 38996 0 1 12562
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_13
timestamp 1624127230
transform 1 0 37670 0 1 12562
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_26
timestamp 1624127230
transform 1 0 40996 0 1 12562
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_29
timestamp 1624127230
transform 1 0 43196 0 1 12562
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_31
timestamp 1624127230
transform 1 0 45196 0 1 12562
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_14
timestamp 1624127230
transform -1 0 46686 0 1 12564
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_14
timestamp 1624127230
transform -1 0 38551 0 1 14176
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_8
timestamp 1624127230
transform -1 0 38529 0 1 14948
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_9
timestamp 1624127230
transform 1 0 37648 0 1 16566
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_21
timestamp 1624127230
transform 1 0 39126 0 1 16580
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_14
timestamp 1624127230
transform 1 0 41034 0 1 14176
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_4
timestamp 1624127230
transform 1 0 41012 0 1 14948
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_20
timestamp 1624127230
transform 1 0 41126 0 1 16580
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_15
timestamp 1624127230
transform -1 0 43322 0 1 14178
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_15
timestamp 1624127230
transform 1 0 45805 0 1 14178
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_9
timestamp 1624127230
transform 1 0 43248 0 1 14948
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_18
timestamp 1624127230
transform 1 0 43326 0 1 16580
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_8
timestamp 1624127230
transform -1 0 45356 0 1 14952
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_19
timestamp 1624127230
transform 1 0 45326 0 1 16580
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_6
timestamp 1624127230
transform -1 0 47678 0 1 14952
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_14
timestamp 1624127230
transform 1 0 47526 0 1 16580
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_10
timestamp 1624127230
transform 1 0 50161 0 1 14952
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_15
timestamp 1624127230
transform 1 0 49526 0 1 16580
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_11
timestamp 1624127230
transform -1 0 51042 0 1 16570
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_8
timestamp 1624127230
transform 1 0 37648 0 1 18670
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_9
timestamp 1624127230
transform -1 0 38529 0 1 20284
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_22
timestamp 1624127230
transform 1 0 39126 0 1 18680
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_23
timestamp 1624127230
transform 1 0 41126 0 1 18680
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_5
timestamp 1624127230
transform 1 0 41012 0 1 20284
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_17
timestamp 1624127230
transform 1 0 43326 0 1 18680
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_16
timestamp 1624127230
transform 1 0 45326 0 1 18680
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_11
timestamp 1624127230
transform 1 0 43248 0 -1 20291
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_10
timestamp 1624127230
transform -1 0 45356 0 -1 20287
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_13
timestamp 1624127230
transform 1 0 47526 0 1 18680
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_JJFNVY  sky130_fd_pr__cap_mim_m3_1_JJFNVY_7
timestamp 1624127230
transform -1 0 47678 0 1 20288
box -950 -300 818 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_12
timestamp 1624127230
transform 1 0 49526 0 1 18680
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_11
timestamp 1624127230
transform 1 0 50161 0 1 20288
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_10
timestamp 1624127230
transform -1 0 51042 0 1 18674
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_3
timestamp 1624127230
transform 1 0 37654 0 1 22616
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_2
timestamp 1624127230
transform -1 0 38535 0 1 21198
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_2
timestamp 1624127230
transform 1 0 37654 0 1 24720
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_2
timestamp 1624127230
transform 1 0 39016 0 1 22614
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_1
timestamp 1624127230
transform 1 0 39016 0 1 24714
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_3
timestamp 1624127230
transform 1 0 41016 0 1 22614
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_3
timestamp 1624127230
transform 1 0 41418 0 1 21198
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_RR5544  sky130_fd_pr__cap_mim_m3_1_RR5544_0
timestamp 1624127230
transform 1 0 41016 0 1 24714
box -950 -900 838 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_1
timestamp 1624127230
transform 1 0 42654 0 1 22616
box -350 -900 244 900
use sky130_fd_pr__cap_mim_m3_1_GJFTVY  sky130_fd_pr__cap_mim_m3_1_GJFTVY_0
timestamp 1624127230
transform 1 0 42654 0 1 24720
box -350 -900 244 900
use txgate  txgate_2
timestamp 1624127230
transform 1 0 -26957 0 1 -35578
box 74185 57360 76542 59116
use txgate  txgate_3
timestamp 1624127230
transform 1 0 -26957 0 1 -33578
box 74185 57360 76542 59116
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_1
timestamp 1624127230
transform -1 0 38535 0 1 26134
box -1350 -300 1232 300
use sky130_fd_pr__cap_mim_m3_1_ZE2L9R  sky130_fd_pr__cap_mim_m3_1_ZE2L9R_0
timestamp 1624127230
transform 1 0 41418 0 1 26134
box -1350 -300 1232 300
use diff_fold_casc_ota  diff_fold_casc_ota_1
timestamp 1624135731
transform 1 0 64950 0 1 26540
box -12400 -27258 25000 1800
<< labels >>
flabel metal3 -9338 5730 -9298 5762 1 FreeSans 480 0 0 0 vhpf
flabel metal3 -9718 1424 -9700 1438 1 FreeSans 480 0 0 0 vincm
flabel metal4 -9700 5602 -9690 5614 1 FreeSans 480 0 0 0 vip1
flabel metal4 -9752 1570 -9732 1586 1 FreeSans 480 0 0 0 vim1
flabel metal3 -9740 8648 -9714 8668 1 FreeSans 480 0 0 0 vim1
flabel metal4 -9698 8802 -9654 8828 1 FreeSans 480 0 0 0 vop1
flabel metal3 -9694 12970 -9674 12986 1 FreeSans 480 0 0 0 vip1
flabel metal4 -9704 12846 -9684 12872 1 FreeSans 480 0 0 0 vom1
flabel metal4 -5616 -342 -5562 -296 1 FreeSans 480 0 0 0 VSS
flabel metal3 39912 1728 39926 1742 1 FreeSans 480 0 0 0 vop1
flabel metal4 39914 1890 39924 1898 1 FreeSans 480 0 0 0 venp1
flabel metal3 39900 6058 39910 6070 1 FreeSans 480 0 0 0 vom1
flabel metal4 39912 5932 39922 5950 1 FreeSans 480 0 0 0 venm1
flabel metal3 39924 13672 39940 13684 1 FreeSans 480 0 0 0 vom1
flabel metal3 39848 9318 39866 9340 1 FreeSans 480 0 0 0 vop1
flabel metal4 39872 9472 39892 9486 1 FreeSans 480 0 0 0 vim2
flabel metal4 39942 13524 39962 13540 1 FreeSans 480 0 0 0 vip2
flabel metal3 40076 15448 40096 15460 1 FreeSans 480 0 0 0 vim2
flabel metal4 40082 15590 40102 15606 1 FreeSans 480 0 0 0 venp2
flabel metal3 40106 19776 40122 19788 1 FreeSans 480 0 0 0 vip2
flabel metal4 40024 19636 40048 19656 1 FreeSans 480 0 0 0 venm2
flabel metal4 40068 25698 40084 25712 1 FreeSans 480 0 0 0 vop
flabel metal3 40216 23534 40238 23550 1 FreeSans 480 0 0 0 vim2
flabel metal4 39646 23652 39664 23674 1 FreeSans 480 0 0 0 vip2
flabel metal4 41908 23258 41930 23278 1 FreeSans 480 0 0 0 vom
flabel metal4 49508 27900 49618 28008 1 FreeSans 480 0 0 0 VDD
flabel metal2 50956 4528 50982 4554 1 FreeSans 480 0 0 0 gain_ctrl_0
flabel metal2 49538 23440 49558 23458 1 FreeSans 480 0 0 0 gain_ctrl_1
flabel metal4 36296 7672 36328 7702 1 FreeSans 480 0 0 0 vocm
flabel metal1 3968 4954 3982 4962 1 FreeSans 480 0 0 0 ibiasn1
flabel metal1 57962 4966 57978 4972 1 FreeSans 480 0 0 0 ibiasn2
flabel metal1 -7768 15456 -7762 15460 1 FreeSans 480 0 0 0 rst_n
flabel metal1 -8136 15450 -8128 15458 1 FreeSans 480 0 0 0 rst
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< error_p >>
rect -29 137 29 143
rect -29 103 -17 137
rect -29 97 29 103
rect -29 -103 29 -97
rect -29 -137 -17 -103
rect -29 -143 29 -137
<< pwell >>
rect -211 -275 211 275
rect -191 -279 211 -275
<< nmos >>
rect -15 -65 15 65
<< ndiff >>
rect -73 53 -15 65
rect -73 -53 -61 53
rect -27 -53 -15 53
rect -73 -65 -15 -53
rect 15 53 73 65
rect 15 -53 27 53
rect 61 -53 73 53
rect 15 -65 73 -53
<< ndiffc >>
rect -61 -53 -27 53
rect 27 -53 61 53
<< psubdiff >>
rect -175 225 -79 259
rect 79 225 175 259
rect -175 86 -141 225
rect 141 86 175 225
rect -175 -239 -141 -86
rect 141 -239 175 -86
rect -175 -273 -79 -239
rect 79 -273 175 -239
<< psubdiffcont >>
rect -79 225 79 259
rect -175 -86 -141 86
rect 141 -86 175 86
rect -79 -273 79 -239
<< poly >>
rect -33 137 33 153
rect -33 103 -17 137
rect 17 103 33 137
rect -33 87 33 103
rect -15 65 15 87
rect -15 -87 15 -65
rect -33 -103 33 -87
rect -33 -137 -17 -103
rect 17 -137 33 -103
rect -33 -153 33 -137
<< polycont >>
rect -17 103 17 137
rect -17 -137 17 -103
<< locali >>
rect -175 225 -79 259
rect 79 225 175 259
rect -175 86 -141 225
rect -33 103 -17 137
rect 17 103 33 137
rect 141 86 175 225
rect -61 53 -27 69
rect -61 -69 -27 -53
rect 27 53 61 69
rect 27 -69 61 -53
rect -175 -239 -141 -86
rect -33 -137 -17 -103
rect 17 -137 33 -103
rect 141 -239 175 -86
rect -175 -273 -79 -239
rect 79 -273 175 -239
<< viali >>
rect -17 103 17 137
rect -61 -53 -27 53
rect 27 -53 61 53
rect -17 -137 17 -103
<< metal1 >>
rect -29 137 29 143
rect -29 103 -17 137
rect 17 103 29 137
rect -29 97 29 103
rect -67 53 -21 65
rect -67 -53 -61 53
rect -27 -53 -21 53
rect -67 -65 -21 -53
rect 21 53 67 65
rect 21 -53 27 53
rect 61 -53 67 53
rect 21 -65 67 -53
rect -29 -103 29 -97
rect -29 -137 -17 -103
rect 17 -137 29 -103
rect -29 -143 29 -137
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string FIXED_BBOX -158 -222 158 222
string parameters w 0.650 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 60 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>

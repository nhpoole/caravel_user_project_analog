magic
tech sky130A
magscale 1 2
timestamp 1624300568
<< nwell >>
rect -3358 -906 2840 2026
rect -3358 -2050 102 -906
rect -3358 -2066 -1014 -2050
rect 76 -2066 102 -2050
<< pwell >>
rect 386 -972 1356 -962
rect 1474 -972 2840 -962
rect 386 -2952 2840 -972
<< psubdiff >>
rect 892 -1476 1054 -1376
rect 2038 -1476 2250 -1376
rect 892 -1538 992 -1476
rect 2150 -1540 2250 -1476
rect 892 -2634 992 -2100
rect 2150 -2634 2250 -2174
rect 892 -2734 1048 -2634
rect 2032 -2734 2250 -2634
<< nsubdiff >>
rect -3322 1890 -3160 1990
rect -120 1890 42 1990
rect -3322 1828 -3222 1890
rect -3322 -1254 -3222 -1192
rect -58 1828 42 1890
rect 380 1890 542 1990
rect 2622 1890 2784 1990
rect 380 1828 480 1890
rect 380 -460 480 -398
rect 2684 1828 2784 1890
rect 2684 -460 2784 -398
rect 380 -560 542 -460
rect 2622 -560 2784 -460
rect -58 -1254 42 -1192
rect -3322 -1354 -3160 -1254
rect -120 -1354 42 -1254
rect -1365 -1415 -7 -1414
rect -1365 -1448 40 -1415
rect -1365 -1449 -1340 -1448
rect -1344 -1450 -1340 -1449
rect 6 -1489 40 -1448
<< psubdiffcont >>
rect 1054 -1476 2038 -1376
rect 892 -2100 992 -1538
rect 2150 -2174 2250 -1540
rect 1048 -2734 2032 -2634
<< nsubdiffcont >>
rect -3160 1890 -120 1990
rect -3322 -1192 -3222 1828
rect -58 -1192 42 1828
rect 542 1890 2622 1990
rect 380 -398 480 1828
rect 2684 -398 2784 1828
rect 542 -560 2622 -460
rect -3160 -1354 -120 -1254
<< poly >>
rect -1092 -1517 -1010 -1507
rect -1092 -1567 -1076 -1517
rect -1026 -1567 -1010 -1517
rect -1092 -1577 -1010 -1567
rect -964 -1517 -882 -1507
rect -964 -1567 -948 -1517
rect -898 -1567 -882 -1517
rect -964 -1577 -882 -1567
rect -836 -1517 -754 -1507
rect -836 -1567 -820 -1517
rect -770 -1567 -754 -1517
rect -836 -1577 -754 -1567
rect -708 -1517 -626 -1507
rect -708 -1567 -692 -1517
rect -642 -1567 -626 -1517
rect -708 -1577 -626 -1567
rect -580 -1517 -498 -1507
rect -580 -1567 -564 -1517
rect -514 -1567 -498 -1517
rect -580 -1577 -498 -1567
rect -452 -1517 -370 -1507
rect -452 -1567 -436 -1517
rect -386 -1567 -370 -1517
rect -452 -1577 -370 -1567
rect -324 -1517 -242 -1507
rect -324 -1567 -308 -1517
rect -258 -1567 -242 -1517
rect -324 -1577 -242 -1567
rect -1086 -1624 -1016 -1577
rect -958 -1624 -888 -1577
rect -830 -1624 -760 -1577
rect -702 -1622 -632 -1577
rect -574 -1623 -504 -1577
rect -446 -1623 -376 -1577
rect -318 -1623 -248 -1577
rect -1214 -1869 -1144 -1824
rect -190 -1869 -120 -1826
rect -1220 -1879 -1138 -1869
rect -1220 -1929 -1204 -1879
rect -1154 -1929 -1138 -1879
rect -1220 -1939 -1138 -1929
rect -196 -1879 -114 -1869
rect -196 -1929 -180 -1879
rect -130 -1929 -114 -1879
rect -196 -1939 -114 -1929
rect 1248 -1542 1308 -1526
rect 1248 -1582 1258 -1542
rect 1298 -1582 1308 -1542
rect 1248 -1644 1308 -1582
rect 1478 -1542 1550 -1532
rect 1478 -1582 1494 -1542
rect 1534 -1582 1550 -1542
rect 1478 -1592 1550 -1582
rect 1596 -1542 1668 -1532
rect 1596 -1582 1612 -1542
rect 1652 -1582 1668 -1542
rect 1596 -1592 1668 -1582
rect 1832 -1542 1904 -1532
rect 1832 -1582 1848 -1542
rect 1888 -1582 1904 -1542
rect 1832 -1592 1904 -1582
rect 1484 -1646 1544 -1592
rect 1602 -1646 1662 -1592
rect 1838 -1644 1898 -1592
rect 1130 -1896 1190 -1848
rect 1064 -1906 1190 -1896
rect 1366 -1898 1426 -1846
rect 1720 -1898 1780 -1846
rect 1956 -1896 2016 -1848
rect 1064 -1946 1080 -1906
rect 1120 -1946 1190 -1906
rect 1064 -1956 1190 -1946
rect 1360 -1908 1432 -1898
rect 1360 -1948 1376 -1908
rect 1416 -1948 1432 -1908
rect 1360 -1958 1432 -1948
rect 1714 -1908 1786 -1898
rect 1714 -1948 1730 -1908
rect 1770 -1948 1786 -1908
rect 1714 -1958 1786 -1948
rect 1956 -1906 2084 -1896
rect 1956 -1946 2028 -1906
rect 2068 -1946 2084 -1906
rect 1956 -1956 2084 -1946
<< polycont >>
rect -1076 -1567 -1026 -1517
rect -948 -1567 -898 -1517
rect -820 -1567 -770 -1517
rect -692 -1567 -642 -1517
rect -564 -1567 -514 -1517
rect -436 -1567 -386 -1517
rect -308 -1567 -258 -1517
rect -1204 -1929 -1154 -1879
rect -180 -1929 -130 -1879
rect 1258 -1582 1298 -1542
rect 1494 -1582 1534 -1542
rect 1612 -1582 1652 -1542
rect 1848 -1582 1888 -1542
rect 1080 -1946 1120 -1906
rect 1376 -1948 1416 -1908
rect 1730 -1948 1770 -1908
rect 2028 -1946 2068 -1906
<< locali >>
rect -3322 1828 -3222 1990
rect -3322 -1354 -3222 -1192
rect -58 1828 42 1990
rect 380 1828 480 1990
rect 380 -560 480 -398
rect 2684 1828 2784 1990
rect 2684 -560 2784 -398
rect 1353 -638 1480 -605
rect 1514 -638 1572 -605
rect 1606 -638 1667 -605
rect 1353 -639 1667 -638
rect 1357 -1150 1572 -1149
rect 1357 -1183 1480 -1150
rect 1514 -1182 1572 -1150
rect 1606 -1182 1715 -1149
rect 1514 -1183 1715 -1182
rect -58 -1354 42 -1192
rect -1347 -1448 -1278 -1414
rect -54 -1415 -12 -1414
rect -54 -1448 40 -1415
rect -1347 -1449 -1340 -1448
rect -1344 -1450 -1340 -1449
rect 6 -1495 40 -1448
rect -1076 -1512 -1026 -1501
rect -948 -1512 -898 -1501
rect -820 -1512 -770 -1501
rect -692 -1507 -642 -1501
rect -564 -1507 -514 -1501
rect -436 -1507 -386 -1501
rect -308 -1507 -258 -1501
rect -702 -1512 -189 -1507
rect -1212 -1517 -189 -1512
rect -1212 -1567 -1076 -1517
rect -1026 -1567 -948 -1517
rect -898 -1567 -820 -1517
rect -770 -1567 -692 -1517
rect -642 -1567 -564 -1517
rect -514 -1567 -436 -1517
rect -386 -1567 -308 -1517
rect -258 -1567 -189 -1517
rect -1212 -1572 -189 -1567
rect -1076 -1583 -1026 -1572
rect -948 -1583 -898 -1572
rect -820 -1583 -770 -1572
rect -702 -1577 -189 -1572
rect -692 -1583 -642 -1577
rect -564 -1583 -514 -1577
rect -436 -1583 -386 -1577
rect -308 -1583 -258 -1577
rect -1277 -1862 -1207 -1785
rect -125 -1862 -55 -1791
rect -1277 -1863 -1188 -1862
rect -132 -1863 -130 -1862
rect -1204 -1869 -1154 -1863
rect -180 -1869 -130 -1863
rect -1204 -1879 -1144 -1869
rect -1154 -1929 -1144 -1879
rect -1204 -1936 -1144 -1929
rect -1277 -1939 -1144 -1936
rect -190 -1879 -130 -1869
rect -190 -1929 -180 -1879
rect -190 -1937 -130 -1929
rect -190 -1939 -55 -1937
rect -1204 -1945 -1154 -1939
rect -180 -1945 -130 -1939
rect 892 -1517 992 -1376
rect 2150 -1516 2250 -1376
rect 1494 -1532 1652 -1526
rect 1848 -1532 1888 -1526
rect 1484 -1542 1662 -1532
rect 1242 -1582 1248 -1542
rect 1308 -1582 1314 -1542
rect 1484 -1582 1494 -1542
rect 1534 -1582 1612 -1542
rect 1652 -1582 1662 -1542
rect 1484 -1592 1662 -1582
rect 1494 -1598 1652 -1592
rect 1848 -1598 1888 -1592
rect 1542 -1682 1602 -1598
rect 1080 -1896 1120 -1890
rect 1376 -1898 1416 -1892
rect 1730 -1898 1770 -1892
rect 2028 -1896 2068 -1890
rect 1366 -1904 1500 -1898
rect 1366 -1908 1446 -1904
rect 1366 -1948 1376 -1908
rect 1416 -1948 1446 -1908
rect 1366 -1952 1446 -1948
rect 1494 -1952 1500 -1904
rect 1080 -1962 1120 -1956
rect 1366 -1958 1500 -1952
rect 1664 -1904 1780 -1898
rect 1664 -1952 1666 -1904
rect 1714 -1908 1780 -1904
rect 1714 -1948 1730 -1908
rect 1770 -1948 1780 -1908
rect 1714 -1952 1780 -1948
rect 1664 -1958 1780 -1952
rect 1376 -1964 1416 -1958
rect 1730 -1964 1770 -1958
rect 2028 -1962 2068 -1956
rect 892 -2734 992 -2593
rect 2150 -2734 2250 -2593
<< viali >>
rect -3222 1890 -3160 1990
rect -3160 1890 -120 1990
rect -120 1890 -58 1990
rect -3322 -1117 -3222 1753
rect -58 -1117 42 1753
rect 480 1890 542 1990
rect 542 1890 2622 1990
rect 2622 1890 2684 1990
rect 380 -368 480 1798
rect 2688 1564 2784 1798
rect 2684 -368 2784 1564
rect 480 -560 542 -460
rect 542 -560 2622 -460
rect 2622 -560 2684 -460
rect 1480 -638 1514 -604
rect 1572 -638 1606 -604
rect 692 -950 740 -902
rect 804 -950 852 -902
rect 964 -950 1012 -902
rect 1072 -950 1120 -902
rect 1204 -950 1252 -902
rect 1378 -950 1426 -902
rect 1674 -950 1708 -916
rect 1852 -952 1900 -904
rect 1966 -952 2014 -904
rect 2082 -950 2130 -902
rect 2242 -950 2290 -902
rect 2354 -950 2402 -902
rect 1384 -1068 1432 -1020
rect 1664 -1068 1712 -1020
rect 1480 -1184 1514 -1150
rect 1572 -1182 1606 -1148
rect -3222 -1354 -3160 -1254
rect -3160 -1354 -120 -1254
rect -120 -1354 -58 -1254
rect -1278 -1448 -54 -1414
rect -1374 -1952 -1340 -1484
rect -1272 -1572 -1212 -1512
rect -189 -1577 -119 -1507
rect -1277 -1936 -1204 -1863
rect -130 -1937 -55 -1862
rect 6 -1952 40 -1506
rect 992 -1476 1054 -1376
rect 1054 -1476 2038 -1376
rect 2038 -1476 2150 -1376
rect 892 -1538 992 -1517
rect 424 -1948 458 -1654
rect 770 -1948 804 -1654
rect -1280 -2030 -56 -1996
rect 892 -2100 992 -1538
rect 1248 -1542 1308 -1532
rect 1248 -1582 1258 -1542
rect 1258 -1582 1298 -1542
rect 1298 -1582 1308 -1542
rect 1248 -1592 1308 -1582
rect 1838 -1542 1898 -1532
rect 1838 -1582 1848 -1542
rect 1848 -1582 1888 -1542
rect 1888 -1582 1898 -1542
rect 1838 -1592 1898 -1582
rect 2150 -1540 2250 -1516
rect 1070 -1906 1130 -1896
rect 1070 -1946 1080 -1906
rect 1080 -1946 1120 -1906
rect 1120 -1946 1130 -1906
rect 1070 -1956 1130 -1946
rect 1446 -1952 1494 -1904
rect 1666 -1952 1714 -1904
rect 2018 -1906 2078 -1896
rect 2018 -1946 2028 -1906
rect 2028 -1946 2068 -1906
rect 2068 -1946 2078 -1906
rect 2018 -1956 2078 -1946
rect 892 -2593 992 -2100
rect 2150 -2174 2250 -1540
rect 2328 -1948 2362 -1654
rect 2674 -1948 2708 -1654
rect 2150 -2593 2250 -2174
rect 992 -2734 1048 -2634
rect 1048 -2734 2032 -2634
rect 2032 -2734 2150 -2634
<< metal1 >>
rect -3328 1990 48 1996
rect -3328 1890 -3222 1990
rect -58 1890 48 1990
rect -3328 1884 48 1890
rect -3328 1753 -3216 1884
rect -3328 -1117 -3322 1753
rect -3222 1584 -3216 1753
rect -348 1584 -330 1884
rect -3222 1564 -330 1584
rect -64 1753 48 1884
rect -3222 -1117 -3216 1564
rect -3166 710 -3106 1564
rect -2134 1242 -2074 1564
rect -1220 1250 -1160 1564
rect -3048 836 -2988 1122
rect -2820 836 -2760 1042
rect -2590 836 -2530 1144
rect -2364 953 -2304 1043
rect -1908 953 -1848 1044
rect -1676 953 -1616 1136
rect -1450 953 -1390 1040
rect -986 953 -926 1042
rect -2364 893 -926 953
rect -762 836 -702 1137
rect -530 836 -470 1044
rect -304 836 -244 1140
rect -3048 776 -244 836
rect -3166 650 -2802 710
rect -3104 536 -3098 596
rect -3038 536 -3032 596
rect -3098 -992 -3038 536
rect -2990 378 -2930 650
rect -2862 452 -2802 650
rect -2986 -192 -2926 50
rect -2862 -192 -2802 -38
rect -2986 -252 -2802 -192
rect -2986 -500 -2926 -252
rect -2862 -404 -2802 -252
rect -2730 -256 -2670 38
rect -2600 -136 -2540 -41
rect -2606 -196 -2600 -136
rect -2540 -196 -2534 -136
rect -2736 -316 -2730 -256
rect -2670 -316 -2664 -256
rect -2476 -528 -2416 776
rect -2220 654 -2214 714
rect -2154 654 -2148 714
rect -2350 536 -2344 596
rect -2284 536 -2278 596
rect -2344 460 -2284 536
rect -2214 336 -2154 654
rect -2092 536 -2086 596
rect -2026 536 -2020 596
rect -2086 460 -2026 536
rect -2352 -196 -2346 -136
rect -2286 -196 -2280 -136
rect -2092 -196 -2086 -136
rect -2026 -196 -2020 -136
rect -2346 -408 -2286 -196
rect -2222 -316 -2216 -256
rect -2156 -316 -2150 -256
rect -2216 -502 -2156 -316
rect -2086 -406 -2026 -196
rect -1958 -516 -1898 776
rect -1828 -136 -1768 -38
rect -1834 -196 -1828 -136
rect -1768 -196 -1762 -136
rect -1700 -256 -1640 60
rect -1570 -136 -1510 -42
rect -1576 -196 -1570 -136
rect -1510 -196 -1504 -136
rect -1706 -316 -1700 -256
rect -1640 -316 -1634 -256
rect -1442 -526 -1382 776
rect -1190 654 -1184 714
rect -1124 654 -1118 714
rect -1318 536 -1312 596
rect -1252 536 -1246 596
rect -1312 454 -1252 536
rect -1184 364 -1124 654
rect -1058 536 -1052 596
rect -992 536 -986 596
rect -1052 456 -992 536
rect -1318 -196 -1312 -136
rect -1252 -196 -1246 -136
rect -1060 -196 -1054 -136
rect -994 -196 -988 -136
rect -1312 -404 -1252 -196
rect -1190 -316 -1184 -256
rect -1124 -316 -1118 -256
rect -1184 -516 -1124 -316
rect -1054 -406 -994 -196
rect -928 -526 -868 776
rect -298 654 -292 714
rect -232 654 -226 714
rect -538 536 -474 596
rect -414 536 -350 596
rect -538 454 -478 536
rect -410 352 -350 536
rect -796 -136 -736 -42
rect -802 -196 -796 -136
rect -736 -196 -730 -136
rect -672 -256 -612 84
rect -538 -198 -478 -42
rect -410 -198 -350 64
rect -678 -316 -672 -256
rect -612 -316 -606 -256
rect -538 -258 -350 -198
rect -538 -404 -478 -258
rect -410 -504 -350 -258
rect -2990 -988 -2930 -792
rect -2860 -988 -2800 -900
rect -3104 -1052 -3098 -992
rect -3038 -1052 -3032 -992
rect -2990 -1048 -2800 -988
rect -2730 -1026 -2670 -810
rect -2604 -992 -2544 -901
rect -1828 -992 -1768 -902
rect -2732 -1108 -2670 -1026
rect -2610 -1052 -2604 -992
rect -2544 -1052 -2538 -992
rect -1834 -1052 -1828 -992
rect -1768 -1052 -1762 -992
rect -3328 -1248 -3216 -1117
rect -2738 -1168 -2732 -1108
rect -2672 -1168 -2666 -1108
rect -1700 -1110 -1640 -792
rect -1572 -992 -1512 -902
rect -800 -992 -740 -898
rect -1578 -1052 -1572 -992
rect -1512 -1052 -1506 -992
rect -806 -1052 -800 -992
rect -740 -1052 -734 -992
rect -1700 -1176 -1640 -1170
rect -670 -1110 -610 -798
rect -538 -990 -478 -904
rect -412 -990 -352 -800
rect -538 -1050 -352 -990
rect -670 -1176 -610 -1170
rect -292 -1110 -232 654
rect -292 -1176 -232 -1170
rect -64 -1117 -58 1753
rect 42 -1117 48 1753
rect 374 1990 2790 1996
rect 374 1890 480 1990
rect 2684 1890 2790 1990
rect 374 1884 2790 1890
rect 374 1798 486 1884
rect 248 366 254 426
rect 314 366 320 426
rect 102 -316 108 -256
rect 168 -316 174 -256
rect -64 -1248 48 -1117
rect -3328 -1254 48 -1248
rect -3328 -1354 -3222 -1254
rect -58 -1354 48 -1254
rect -3328 -1360 48 -1354
rect -1570 -1458 -1564 -1398
rect -1504 -1458 -1498 -1398
rect -1388 -1414 48 -1360
rect -1388 -1448 -1278 -1414
rect -54 -1448 48 -1414
rect -1564 -2076 -1504 -1458
rect -1388 -1462 48 -1448
rect -1388 -1484 -1330 -1462
rect -1388 -1952 -1374 -1484
rect -1340 -1952 -1330 -1484
rect -1278 -1506 -1206 -1500
rect -1284 -1578 -1278 -1506
rect -1218 -1512 -1206 -1506
rect -1212 -1572 -1206 -1512
rect -1218 -1578 -1206 -1572
rect -1278 -1584 -1206 -1578
rect -195 -1501 -113 -1495
rect -195 -1507 -183 -1501
rect -195 -1577 -189 -1507
rect -195 -1583 -183 -1577
rect -113 -1583 -107 -1501
rect -10 -1506 48 -1462
rect -195 -1589 -113 -1583
rect -1276 -1857 -1203 -1786
rect -1152 -1826 -1146 -1766
rect -1086 -1826 -1080 -1766
rect -1289 -1863 -1192 -1857
rect -1289 -1936 -1277 -1863
rect -1204 -1936 -1192 -1863
rect -1016 -1874 -956 -1732
rect -896 -1816 -890 -1756
rect -830 -1816 -824 -1756
rect -762 -1874 -702 -1788
rect -638 -1806 -632 -1746
rect -572 -1806 -566 -1746
rect -506 -1874 -446 -1774
rect -386 -1808 -380 -1748
rect -320 -1808 -314 -1748
rect -252 -1806 -246 -1746
rect -186 -1806 -180 -1746
rect -250 -1874 -190 -1806
rect -129 -1856 -54 -1759
rect -1016 -1934 -190 -1874
rect -142 -1862 -43 -1856
rect -1289 -1942 -1192 -1936
rect -142 -1937 -130 -1862
rect -55 -1937 -43 -1862
rect -1388 -1979 -1330 -1952
rect -1276 -1979 -1203 -1942
rect -142 -1943 -43 -1937
rect -129 -1979 -54 -1943
rect -10 -1952 6 -1506
rect 40 -1952 48 -1506
rect -10 -1979 48 -1952
rect -1388 -1996 48 -1979
rect -1388 -2030 -1280 -1996
rect -56 -2030 48 -1996
rect -1388 -2038 48 -2030
rect -380 -2076 -320 -2070
rect -1564 -2078 -890 -2076
rect -1564 -2136 -1146 -2078
rect -1152 -2138 -1146 -2136
rect -1086 -2136 -890 -2078
rect -830 -2136 -632 -2076
rect -572 -2136 -380 -2076
rect -1086 -2138 -1080 -2136
rect -380 -2142 -320 -2136
rect 108 -2096 168 -316
rect 254 -896 314 366
rect 374 -368 380 1798
rect 480 -368 486 1798
rect 1038 1584 1056 1884
rect 2676 1798 2790 1884
rect 2676 1584 2688 1798
rect 1038 1564 2688 1584
rect 1090 1414 1150 1564
rect 578 1354 1150 1414
rect 578 1024 638 1354
rect 708 1146 768 1354
rect 834 1244 840 1304
rect 900 1244 906 1304
rect 840 1038 900 1244
rect 374 -454 486 -368
rect 574 492 634 850
rect 708 492 768 644
rect 574 432 768 492
rect 574 -312 634 432
rect 708 278 768 432
rect 964 426 1024 644
rect 834 366 840 426
rect 900 366 906 426
rect 958 366 964 426
rect 1024 366 1030 426
rect 840 64 900 366
rect 1090 150 1150 1354
rect 1220 1244 1226 1304
rect 1286 1244 1292 1304
rect 1478 1244 1484 1304
rect 1544 1244 1550 1304
rect 1226 1138 1286 1244
rect 1484 1134 1544 1244
rect 1354 426 1414 746
rect 1220 366 1226 426
rect 1286 366 1292 426
rect 1348 366 1354 426
rect 1414 366 1420 426
rect 1474 366 1480 426
rect 1540 366 1546 426
rect 1226 276 1286 366
rect 1480 276 1540 366
rect 1606 154 1666 1564
rect 1862 1244 1868 1304
rect 1928 1244 1934 1304
rect 1868 1046 1928 1244
rect 1738 426 1798 648
rect 1996 494 2056 645
rect 2124 498 2184 1564
rect 2260 498 2320 640
rect 2386 498 2446 1564
rect 2502 1244 2508 1304
rect 2568 1244 2574 1304
rect 1990 434 1996 494
rect 2056 434 2062 494
rect 2124 438 2446 498
rect 1732 366 1738 426
rect 1798 366 1804 426
rect 1862 366 1868 426
rect 1928 366 1934 426
rect 1868 172 1928 366
rect 1996 276 2056 434
rect 2124 172 2184 438
rect 2260 284 2320 438
rect 2386 176 2446 438
rect 712 -312 772 -218
rect 574 -372 772 -312
rect 960 -328 1020 -217
rect 1350 -328 1410 -112
rect 1738 -328 1798 -218
rect 2508 -328 2568 1244
rect 954 -388 960 -328
rect 1020 -388 1026 -328
rect 1344 -388 1350 -328
rect 1410 -388 1416 -328
rect 1732 -388 1738 -328
rect 1798 -388 1804 -328
rect 2502 -388 2508 -328
rect 2568 -388 2574 -328
rect 2678 -368 2684 1564
rect 2784 -368 2790 1798
rect 2678 -454 2790 -368
rect 374 -460 2790 -454
rect 374 -560 480 -460
rect 2684 -560 2790 -460
rect 374 -566 2790 -560
rect 626 -604 2470 -566
rect 626 -638 1480 -604
rect 1514 -638 1572 -604
rect 1606 -638 2470 -604
rect 626 -652 2470 -638
rect 1418 -670 1658 -652
rect 2772 -680 2778 -620
rect 2838 -680 2844 -620
rect 798 -896 858 -890
rect 958 -896 1018 -890
rect 254 -902 752 -896
rect 254 -950 692 -902
rect 740 -950 752 -902
rect 254 -956 752 -950
rect 798 -902 1018 -896
rect 798 -950 804 -902
rect 852 -950 964 -902
rect 1012 -950 1018 -902
rect 798 -956 1018 -950
rect 1060 -902 1264 -896
rect 1060 -950 1072 -902
rect 1120 -950 1204 -902
rect 1252 -950 1264 -902
rect 1060 -956 1264 -950
rect 1366 -902 1612 -896
rect 1366 -950 1378 -902
rect 1426 -950 1612 -902
rect 1846 -898 1906 -892
rect 1960 -898 2020 -892
rect 2076 -896 2136 -890
rect 2236 -896 2296 -890
rect 1846 -904 2028 -898
rect 1366 -956 1612 -950
rect 254 -1988 314 -956
rect 798 -962 858 -956
rect 958 -962 1018 -956
rect 1378 -1014 1438 -1008
rect 1552 -1014 1612 -956
rect 1652 -964 1658 -904
rect 1718 -964 1724 -904
rect 1846 -952 1852 -904
rect 1900 -952 1966 -904
rect 2014 -952 2028 -904
rect 1846 -958 2028 -952
rect 2076 -902 2296 -896
rect 2076 -950 2082 -902
rect 2130 -950 2242 -902
rect 2290 -950 2296 -902
rect 2076 -956 2296 -950
rect 1846 -964 1906 -958
rect 1960 -964 2020 -958
rect 2076 -962 2136 -956
rect 2236 -962 2296 -956
rect 2348 -896 2408 -890
rect 2778 -896 2838 -680
rect 2348 -902 2838 -896
rect 2348 -950 2354 -902
rect 2402 -950 2838 -902
rect 2348 -956 2838 -950
rect 2348 -962 2408 -956
rect 1658 -1014 1718 -1008
rect 1372 -1074 1378 -1014
rect 1438 -1074 1444 -1014
rect 1552 -1020 1718 -1014
rect 1552 -1068 1664 -1020
rect 1712 -1068 1718 -1020
rect 1552 -1074 1718 -1068
rect 1378 -1080 1438 -1074
rect 1658 -1080 1718 -1074
rect 1446 -1120 1686 -1118
rect 972 -1148 2110 -1120
rect 972 -1150 1572 -1148
rect 972 -1184 1480 -1150
rect 1514 -1182 1572 -1150
rect 1606 -1182 2110 -1148
rect 1514 -1184 2110 -1182
rect 972 -1202 2110 -1184
rect 886 -1376 2256 -1202
rect 886 -1476 992 -1376
rect 2150 -1476 2256 -1376
rect 886 -1482 2256 -1476
rect 886 -1517 998 -1482
rect 412 -1654 472 -1640
rect 412 -1948 424 -1654
rect 458 -1948 472 -1654
rect 558 -1702 564 -1602
rect 664 -1702 670 -1602
rect 756 -1654 820 -1642
rect 248 -2048 254 -1988
rect 314 -2048 320 -1988
rect 108 -2162 168 -2156
rect 412 -2282 472 -1948
rect 526 -1988 586 -1764
rect 642 -1794 702 -1734
rect 642 -1926 704 -1794
rect 642 -1988 702 -1926
rect 756 -1948 770 -1654
rect 804 -1948 820 -1654
rect 520 -2048 526 -1988
rect 586 -2048 592 -1988
rect 636 -2048 642 -1988
rect 702 -2048 708 -1988
rect 756 -2282 820 -1948
rect 886 -2282 892 -1517
rect 322 -2308 892 -2282
rect 992 -2280 998 -1517
rect 2144 -1516 2256 -1482
rect 1130 -1532 1190 -1526
rect 1242 -1532 1314 -1520
rect 1832 -1532 1904 -1520
rect 1190 -1592 1248 -1532
rect 1308 -1592 1838 -1532
rect 1898 -1592 1904 -1532
rect 1130 -1598 1190 -1592
rect 1242 -1604 1314 -1592
rect 1424 -1680 1484 -1592
rect 1662 -1672 1722 -1592
rect 1832 -1604 1904 -1592
rect 1070 -1884 1130 -1814
rect 1064 -1896 1136 -1884
rect 1064 -1956 1070 -1896
rect 1130 -1956 1136 -1896
rect 1064 -1968 1136 -1956
rect 1070 -2280 1130 -1968
rect 1188 -2098 1248 -1814
rect 1182 -2158 1188 -2098
rect 1248 -2158 1254 -2098
rect 1310 -2280 1370 -1808
rect 1440 -1898 1500 -1892
rect 1434 -1958 1440 -1898
rect 1500 -1958 1506 -1898
rect 1440 -1964 1500 -1958
rect 1542 -2280 1602 -1822
rect 1660 -1898 1720 -1892
rect 1654 -1958 1660 -1898
rect 1720 -1958 1726 -1898
rect 1660 -1964 1720 -1958
rect 1778 -2280 1838 -1810
rect 1896 -2098 1956 -1810
rect 2018 -1884 2078 -1792
rect 2012 -1896 2084 -1884
rect 2012 -1956 2018 -1896
rect 2078 -1956 2084 -1896
rect 2012 -1968 2084 -1956
rect 1890 -2158 1896 -2098
rect 1956 -2158 1962 -2098
rect 2018 -2280 2078 -1968
rect 2144 -2280 2150 -1516
rect 992 -2308 2150 -2280
rect 2250 -2280 2256 -1516
rect 2316 -1654 2376 -1642
rect 2316 -1948 2328 -1654
rect 2362 -1948 2376 -1654
rect 2462 -1704 2468 -1604
rect 2568 -1704 2574 -1604
rect 2662 -1654 2722 -1644
rect 2316 -2280 2376 -1948
rect 2426 -2098 2486 -1884
rect 2546 -1998 2606 -1878
rect 2662 -1948 2674 -1654
rect 2708 -1948 2722 -1654
rect 2540 -2058 2546 -1998
rect 2606 -2058 2612 -1998
rect 2420 -2158 2426 -2098
rect 2486 -2158 2492 -2098
rect 2662 -2280 2722 -1948
rect 2778 -1998 2838 -956
rect 2772 -2058 2778 -1998
rect 2838 -2058 2844 -1998
rect 2250 -2308 2810 -2280
rect 322 -2614 346 -2308
rect 2790 -2614 2810 -2308
rect 322 -2632 2810 -2614
rect 886 -2634 2256 -2632
rect 886 -2734 992 -2634
rect 2150 -2734 2256 -2634
rect 886 -2740 2256 -2734
<< via1 >>
rect -3216 1584 -348 1884
rect -3098 536 -3038 596
rect -2600 -196 -2540 -136
rect -2730 -316 -2670 -256
rect -2214 654 -2154 714
rect -2344 536 -2284 596
rect -2086 536 -2026 596
rect -2346 -196 -2286 -136
rect -2086 -196 -2026 -136
rect -2216 -316 -2156 -256
rect -1828 -196 -1768 -136
rect -1570 -196 -1510 -136
rect -1700 -316 -1640 -256
rect -1184 654 -1124 714
rect -1312 536 -1252 596
rect -1052 536 -992 596
rect -1312 -196 -1252 -136
rect -1054 -196 -994 -136
rect -1184 -316 -1124 -256
rect -292 654 -232 714
rect -474 536 -414 596
rect -796 -196 -736 -136
rect -672 -316 -612 -256
rect -3098 -1052 -3038 -992
rect -2604 -1052 -2544 -992
rect -1828 -1052 -1768 -992
rect -2732 -1168 -2672 -1108
rect -1572 -1052 -1512 -992
rect -800 -1052 -740 -992
rect -1700 -1170 -1640 -1110
rect -670 -1170 -610 -1110
rect -292 -1170 -232 -1110
rect 254 366 314 426
rect 108 -316 168 -256
rect -1564 -1458 -1504 -1398
rect -1278 -1512 -1218 -1506
rect -1278 -1572 -1272 -1512
rect -1272 -1572 -1218 -1512
rect -1278 -1578 -1218 -1572
rect -183 -1507 -113 -1501
rect -183 -1577 -119 -1507
rect -119 -1577 -113 -1507
rect -183 -1583 -113 -1577
rect -1146 -1826 -1086 -1766
rect -890 -1816 -830 -1756
rect -632 -1806 -572 -1746
rect -380 -1808 -320 -1748
rect -246 -1806 -186 -1746
rect -1146 -2138 -1086 -2078
rect -890 -2136 -830 -2076
rect -632 -2136 -572 -2076
rect -380 -2136 -320 -2076
rect 1056 1584 2676 1884
rect 840 1244 900 1304
rect 840 366 900 426
rect 964 366 1024 426
rect 1226 1244 1286 1304
rect 1484 1244 1544 1304
rect 1226 366 1286 426
rect 1354 366 1414 426
rect 1480 366 1540 426
rect 1868 1244 1928 1304
rect 2508 1244 2568 1304
rect 1996 434 2056 494
rect 1738 366 1798 426
rect 1868 366 1928 426
rect 960 -388 1020 -328
rect 1350 -388 1410 -328
rect 1738 -388 1798 -328
rect 2508 -388 2568 -328
rect 2778 -680 2838 -620
rect 1658 -916 1718 -904
rect 1658 -950 1674 -916
rect 1674 -950 1708 -916
rect 1708 -950 1718 -916
rect 1658 -964 1718 -950
rect 1378 -1020 1438 -1014
rect 1378 -1068 1384 -1020
rect 1384 -1068 1432 -1020
rect 1432 -1068 1438 -1020
rect 1378 -1074 1438 -1068
rect 564 -1702 664 -1602
rect 254 -2048 314 -1988
rect 108 -2156 168 -2096
rect 526 -2048 586 -1988
rect 642 -2048 702 -1988
rect 1130 -1592 1190 -1532
rect 1188 -2158 1248 -2098
rect 1440 -1904 1500 -1898
rect 1440 -1952 1446 -1904
rect 1446 -1952 1494 -1904
rect 1494 -1952 1500 -1904
rect 1440 -1958 1500 -1952
rect 1660 -1904 1720 -1898
rect 1660 -1952 1666 -1904
rect 1666 -1952 1714 -1904
rect 1714 -1952 1720 -1904
rect 1660 -1958 1720 -1952
rect 1896 -2158 1956 -2098
rect 2468 -1704 2568 -1604
rect 2546 -2058 2606 -1998
rect 2426 -2158 2486 -2098
rect 2778 -2058 2838 -1998
rect 346 -2593 892 -2308
rect 892 -2593 992 -2308
rect 992 -2593 2150 -2308
rect 2150 -2593 2250 -2308
rect 2250 -2593 2790 -2308
rect 346 -2614 2790 -2593
<< metal2 >>
rect -3216 1884 -348 1894
rect 1056 1884 2676 1894
rect -348 1584 -112 1650
rect -3216 1574 -112 1584
rect 1056 1574 2676 1584
rect -2214 714 -2154 720
rect -1184 714 -1124 720
rect -292 714 -232 720
rect -2154 654 -1184 714
rect -1124 654 -292 714
rect -2214 648 -2154 654
rect -1184 648 -1124 654
rect -292 648 -232 654
rect -3098 596 -3038 602
rect -2344 596 -2284 602
rect -2086 596 -2026 602
rect -1312 596 -1252 602
rect -1052 596 -992 602
rect -3038 536 -2344 596
rect -2284 536 -2086 596
rect -2026 536 -1312 596
rect -1252 536 -1052 596
rect -3098 530 -3038 536
rect -2344 530 -2284 536
rect -2086 530 -2026 536
rect -1312 530 -1252 536
rect -1052 530 -992 536
rect -474 596 -414 602
rect -172 596 -112 1574
rect 840 1304 900 1310
rect 1226 1304 1286 1310
rect 1484 1304 1544 1310
rect 1868 1304 1928 1310
rect 2508 1304 2568 1310
rect 900 1244 1226 1304
rect 1286 1244 1484 1304
rect 1544 1244 1868 1304
rect 1928 1244 2508 1304
rect 840 1238 900 1244
rect 1226 1238 1286 1244
rect 1484 1238 1544 1244
rect 1868 1238 1928 1244
rect 2508 1238 2568 1244
rect -414 536 -112 596
rect -474 530 -414 536
rect 1996 494 2056 500
rect 1987 434 1996 494
rect 2056 434 2065 494
rect 254 426 314 432
rect 840 426 900 432
rect 964 426 1024 432
rect 1226 426 1286 432
rect 1354 426 1414 432
rect 1480 426 1540 432
rect 1738 426 1798 432
rect 1868 426 1928 432
rect 1996 428 2056 434
rect 314 366 840 426
rect 900 366 964 426
rect 1024 366 1226 426
rect 1286 366 1354 426
rect 1414 366 1480 426
rect 1540 366 1738 426
rect 1798 366 1868 426
rect 254 360 314 366
rect 840 360 900 366
rect 964 360 1024 366
rect 1226 360 1286 366
rect 1354 360 1414 366
rect 1480 360 1540 366
rect 1738 360 1798 366
rect 1868 360 1928 366
rect -2600 -136 -2540 -130
rect -2346 -136 -2286 -130
rect -2086 -136 -2026 -130
rect -1828 -136 -1768 -130
rect -1570 -136 -1510 -130
rect -1312 -136 -1252 -130
rect -1054 -136 -994 -130
rect -796 -136 -736 -130
rect -2540 -196 -2346 -136
rect -2286 -196 -2086 -136
rect -2026 -196 -1828 -136
rect -1768 -196 -1570 -136
rect -1510 -196 -1312 -136
rect -1252 -196 -1054 -136
rect -994 -196 -796 -136
rect -2600 -202 -2540 -196
rect -2346 -202 -2286 -196
rect -2086 -202 -2026 -196
rect -1828 -202 -1768 -196
rect -1570 -202 -1510 -196
rect -1312 -202 -1252 -196
rect -1054 -202 -994 -196
rect -796 -202 -736 -196
rect -2730 -256 -2670 -250
rect -2216 -256 -2156 -250
rect -1700 -256 -1640 -250
rect -1184 -256 -1124 -250
rect -672 -256 -612 -250
rect 108 -256 168 -250
rect -2670 -316 -2216 -256
rect -2156 -316 -1700 -256
rect -1640 -316 -1184 -256
rect -1124 -316 -672 -256
rect -612 -316 108 -256
rect -2730 -322 -2670 -316
rect -2216 -322 -2156 -316
rect -1700 -322 -1640 -316
rect -1184 -322 -1124 -316
rect -672 -322 -612 -316
rect 108 -322 168 -316
rect 960 -328 1020 -322
rect 1350 -328 1410 -322
rect 1738 -328 1798 -322
rect 2508 -328 2568 -322
rect 1020 -388 1350 -328
rect 1410 -388 1738 -328
rect 1798 -388 2508 -328
rect 2568 -388 2838 -328
rect 960 -394 1020 -388
rect 1350 -394 1410 -388
rect 1738 -394 1798 -388
rect 2508 -394 2568 -388
rect 1484 -570 2616 -510
rect 1484 -904 1544 -570
rect 1658 -904 1718 -898
rect 1484 -964 1658 -904
rect -3098 -992 -3038 -986
rect -2604 -992 -2544 -986
rect -1828 -992 -1768 -986
rect -1572 -992 -1512 -986
rect -800 -992 -740 -986
rect -3038 -1052 -2604 -992
rect -2544 -1052 -1828 -992
rect -1768 -1052 -1572 -992
rect -1512 -1052 -800 -992
rect -3098 -1058 -3038 -1052
rect -2604 -1058 -2544 -1052
rect -1828 -1058 -1768 -1052
rect -1572 -1058 -1512 -1052
rect -800 -1058 -740 -1052
rect 1378 -1014 1438 -1008
rect 1484 -1014 1544 -964
rect 1658 -970 1718 -964
rect 2556 -962 2616 -570
rect 2778 -620 2838 -388
rect 2778 -686 2838 -680
rect 1438 -1074 1544 -1014
rect 2556 -1022 2844 -962
rect 1378 -1080 1438 -1074
rect -2732 -1108 -2672 -1102
rect -2672 -1110 586 -1108
rect -2672 -1168 -1700 -1110
rect -2732 -1174 -2672 -1168
rect -1706 -1170 -1700 -1168
rect -1640 -1168 -670 -1110
rect -1640 -1170 -1634 -1168
rect -1564 -1398 -1504 -1168
rect -676 -1170 -670 -1168
rect -610 -1168 -292 -1110
rect -610 -1170 -604 -1168
rect -298 -1170 -292 -1168
rect -232 -1168 586 -1110
rect -232 -1170 -226 -1168
rect 526 -1208 586 -1168
rect 526 -1268 1018 -1208
rect -1564 -1464 -1504 -1458
rect -1278 -1506 -1218 -1500
rect -183 -1501 -113 -1495
rect -1287 -1578 -1278 -1506
rect -1218 -1578 -1209 -1506
rect -1278 -1584 -1218 -1578
rect -192 -1583 -183 -1501
rect -113 -1583 -104 -1501
rect 958 -1532 1018 -1268
rect -183 -1589 -113 -1583
rect 958 -1592 1130 -1532
rect 1190 -1592 1196 -1532
rect 564 -1602 664 -1596
rect 560 -1697 564 -1607
rect 664 -1697 668 -1607
rect 564 -1708 664 -1702
rect -632 -1746 -572 -1740
rect -890 -1756 -830 -1750
rect -1146 -1766 -1086 -1760
rect -1146 -2078 -1086 -1826
rect -1146 -2144 -1086 -2138
rect -890 -2076 -830 -1816
rect -890 -2142 -830 -2136
rect -632 -2076 -572 -1806
rect -380 -1748 -320 -1742
rect -380 -2076 -320 -1808
rect -246 -1746 -186 -1740
rect -386 -2136 -380 -2076
rect -320 -2136 -314 -2076
rect -246 -2098 -186 -1806
rect 254 -1988 314 -1982
rect 526 -1988 586 -1982
rect 642 -1988 702 -1982
rect 958 -1988 1018 -1592
rect 2468 -1604 2568 -1598
rect 2464 -1699 2468 -1609
rect 2568 -1699 2572 -1609
rect 2468 -1710 2568 -1704
rect 1434 -1958 1440 -1898
rect 1500 -1958 1660 -1898
rect 1720 -1958 1726 -1898
rect 314 -2048 526 -1988
rect 636 -2048 642 -1988
rect 702 -2048 1018 -1988
rect 254 -2054 314 -2048
rect 526 -2054 586 -2048
rect 642 -2054 702 -2048
rect 102 -2098 108 -2096
rect -632 -2142 -572 -2136
rect -246 -2156 108 -2098
rect 168 -2098 174 -2096
rect 1188 -2098 1248 -2092
rect 1542 -2098 1602 -1958
rect 2546 -1998 2606 -1992
rect 2778 -1998 2838 -1992
rect 2606 -2058 2778 -1998
rect 2546 -2064 2606 -2058
rect 2778 -2064 2838 -2058
rect 1896 -2098 1956 -2092
rect 2426 -2098 2486 -2092
rect 168 -2156 1188 -2098
rect -246 -2158 1188 -2156
rect 1248 -2158 1896 -2098
rect 1956 -2158 2426 -2098
rect 1188 -2164 1248 -2158
rect 2426 -2164 2486 -2158
rect 346 -2308 2790 -2298
rect 346 -2624 2790 -2614
<< via2 >>
rect -3216 1584 -348 1884
rect 1056 1584 2676 1884
rect 1996 434 2056 494
rect -1278 -1578 -1218 -1506
rect -183 -1583 -113 -1501
rect 569 -1697 659 -1607
rect 2473 -1699 2563 -1609
rect 346 -2614 2790 -2308
<< metal3 >>
rect -3226 1884 -338 1889
rect -3226 1584 -3216 1884
rect -348 1584 -338 1884
rect -3226 1579 -338 1584
rect 1046 1884 2686 1889
rect 1046 1584 1056 1884
rect 2676 1584 2686 1884
rect 1046 1579 2686 1584
rect 1978 499 2078 516
rect 1978 494 1997 499
rect 1978 434 1996 494
rect 1978 429 1997 434
rect 2061 429 2078 499
rect 1978 416 2078 429
rect 2946 -1238 3046 -1232
rect -2188 -1590 -2182 -1490
rect -2082 -1590 -2076 -1490
rect -1298 -1501 -1196 -1492
rect -1298 -1583 -1283 -1501
rect -1219 -1506 -1196 -1501
rect -1218 -1578 -1196 -1506
rect -1219 -1583 -1196 -1578
rect -2182 -2858 -2082 -1590
rect -1298 -1592 -1196 -1583
rect -202 -1496 -96 -1488
rect -202 -1501 -178 -1496
rect -202 -1583 -183 -1501
rect -202 -1588 -178 -1583
rect -108 -1588 -96 -1496
rect -202 -1596 -96 -1588
rect 564 -1603 664 -1602
rect 559 -1701 565 -1603
rect 663 -1701 669 -1603
rect 2468 -1605 2568 -1604
rect 564 -1702 664 -1701
rect 2463 -1703 2469 -1605
rect 2567 -1703 2573 -1605
rect 2468 -1704 2568 -1703
rect 336 -2308 2800 -2303
rect 336 -2614 346 -2308
rect 2790 -2614 2800 -2308
rect 336 -2619 2800 -2614
rect 2946 -2858 3046 -1338
rect -2182 -2958 3046 -2858
<< via3 >>
rect -3216 1584 -348 1884
rect 1056 1584 2676 1884
rect 1997 494 2061 499
rect 1997 434 2056 494
rect 2056 434 2061 494
rect 1997 429 2061 434
rect 2946 -1338 3046 -1238
rect -2182 -1590 -2082 -1490
rect -1283 -1506 -1219 -1501
rect -1283 -1578 -1278 -1506
rect -1278 -1578 -1219 -1506
rect -1283 -1583 -1219 -1578
rect -178 -1501 -108 -1496
rect -178 -1583 -113 -1501
rect -113 -1583 -108 -1501
rect -178 -1588 -108 -1583
rect 565 -1607 663 -1603
rect 565 -1697 569 -1607
rect 569 -1697 659 -1607
rect 659 -1697 663 -1607
rect 565 -1701 663 -1697
rect 2469 -1609 2567 -1605
rect 2469 -1699 2473 -1609
rect 2473 -1699 2563 -1609
rect 2563 -1699 2567 -1609
rect 2469 -1703 2567 -1699
rect 346 -2614 2790 -2308
<< metal4 >>
rect -3400 1884 2890 2278
rect -3400 1584 -3216 1884
rect -348 1584 1056 1884
rect 2676 1584 2890 1884
rect -3400 1478 2890 1584
rect 1976 499 3044 516
rect 1976 429 1997 499
rect 2061 429 3044 499
rect 1976 416 3044 429
rect 2944 -1237 3044 416
rect 2944 -1238 3047 -1237
rect 2944 -1244 2946 -1238
rect 2468 -1338 2946 -1244
rect 3046 -1338 3047 -1238
rect 2468 -1339 3047 -1338
rect 2468 -1344 3044 -1339
rect -2183 -1490 -2081 -1489
rect -2183 -1492 -2182 -1490
rect -2190 -1590 -2182 -1492
rect -2082 -1492 -2081 -1490
rect -2082 -1496 668 -1492
rect -2082 -1501 -178 -1496
rect -2082 -1583 -1283 -1501
rect -1219 -1583 -178 -1501
rect -2082 -1588 -178 -1583
rect -108 -1588 668 -1496
rect -2082 -1590 668 -1588
rect -2190 -1592 668 -1590
rect 564 -1603 668 -1592
rect 564 -1701 565 -1603
rect 663 -1701 668 -1603
rect 564 -1702 668 -1701
rect 568 -1706 668 -1702
rect 2468 -1605 2568 -1344
rect 2468 -1703 2469 -1605
rect 2567 -1703 2568 -1605
rect 2468 -1704 2568 -1703
rect -3400 -2308 2890 -2214
rect -3400 -2614 346 -2308
rect 2790 -2614 2890 -2308
rect -3400 -3014 2890 -2614
use sky130_fd_pr__pfet_01v8_lvt_XJHVCG  sky130_fd_pr__pfet_01v8_lvt_XJHVCG_0
timestamp 1624299007
transform 1 0 -667 0 1 -1724
box -743 -342 743 346
use sky130_fd_pr__nfet_01v8_7DDHNL  sky130_fd_pr__nfet_01v8_7DDHNL_0
timestamp 1624299007
transform 1 0 1573 0 1 -1746
box -501 -126 501 126
use sky130_fd_pr__nfet_01v8_BGQ2FN  sky130_fd_pr__nfet_01v8_BGQ2FN_0
timestamp 1624299007
transform 1 0 614 0 1 -1801
box -226 -279 226 279
use sky130_fd_pr__nfet_01v8_BGQ2FN  sky130_fd_pr__nfet_01v8_BGQ2FN_1
timestamp 1624299007
transform 1 0 2518 0 1 -1801
box -226 -279 226 279
use sky130_fd_pr__pfet_01v8_lvt_JN5RQF  sky130_fd_pr__pfet_01v8_lvt_JN5RQF_1
timestamp 1624299007
transform 1 0 -1670 0 1 -653
box -1355 -300 1355 300
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624299007
transform -1 0 2468 0 1 -1166
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2
timestamp 1624299007
transform -1 0 2192 0 1 -1166
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1624299007
transform 1 0 902 0 1 -1166
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1624299007
transform 1 0 626 0 1 -1166
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_0 ~/PDKS/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624299007
transform 1 0 1178 0 1 -1166
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  sky130_fd_sc_hd__nand2_1_1
timestamp 1624299007
transform -1 0 1916 0 1 -1166
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_lvt_JN5RQF  sky130_fd_pr__pfet_01v8_lvt_JN5RQF_0
timestamp 1624299007
transform 1 0 -1670 0 1 207
box -1355 -300 1355 300
use sky130_fd_pr__pfet_01v8_9JKHSP  sky130_fd_pr__pfet_01v8_9JKHSP_1
timestamp 1624299007
transform 1 0 1512 0 1 30
box -968 -300 968 300
use sky130_fd_pr__pfet_01v8_9JKHSP  sky130_fd_pr__pfet_01v8_9JKHSP_0
timestamp 1624299007
transform 1 0 1512 0 1 890
box -968 -300 968 300
use sky130_fd_pr__pfet_01v8_RCENQY  sky130_fd_pr__pfet_01v8_RCENQY_0
timestamp 1624299007
transform 1 0 -1645 0 1 1190
box -1439 -200 1439 200
<< labels >>
flabel metal4 324 2134 340 2140 1 FreeSans 480 0 0 0 VDD
flabel metal1 -3086 -112 -3072 -100 1 FreeSans 480 0 0 0 vip
flabel metal1 -2316 -232 -2306 -222 1 FreeSans 480 0 0 0 vim
flabel metal1 -276 278 -262 298 1 FreeSans 480 0 0 0 vlatchm
flabel metal1 -2710 -188 -2696 -178 1 FreeSans 480 0 0 0 vlatchp
flabel metal1 -1664 800 -1646 814 1 FreeSans 480 0 0 0 vtailp
flabel metal1 -1746 918 -1726 930 1 FreeSans 480 0 0 0 ibiasp
flabel via1 862 368 878 384 1 FreeSans 480 0 0 0 vcompm
flabel metal1 2526 590 2546 614 1 FreeSans 480 0 0 0 vcompp
flabel metal4 -186 -2534 -160 -2514 1 FreeSans 480 0 0 0 VSS
flabel metal1 1360 -1568 1366 -1562 1 FreeSans 480 0 0 0 vlatchm
flabel metal2 1448 -2134 1456 -2126 1 FreeSans 480 0 0 0 vlatchp
flabel metal1 1156 -934 1162 -928 1 FreeSans 160 0 0 0 vcompm_buf
flabel metal1 900 -934 906 -930 1 FreeSans 160 0 0 0 vcompmb
flabel metal1 1924 -930 1928 -926 1 FreeSans 160 0 0 0 vcompp_buf
flabel metal1 2178 -932 2184 -928 1 FreeSans 160 0 0 0 vcomppb
flabel metal2 2674 -990 2680 -984 1 FreeSans 480 0 0 0 vop
flabel metal1 1606 -1052 1612 -1044 1 FreeSans 480 0 0 0 vom
flabel metal4 -1548 -1552 -1528 -1534 1 FreeSans 480 0 0 0 clk
<< properties >>
string FIXED_BBOX 308 88 2612 2032
<< end >>

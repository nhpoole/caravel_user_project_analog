magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< error_p >>
rect -743 344 743 346
rect -743 248 -731 344
rect -707 308 707 310
rect -707 212 -695 308
<< nwell >>
rect -731 248 743 344
rect -743 -342 743 248
<< pmoslvt >>
rect -547 -100 -477 100
rect -419 -100 -349 100
rect -291 -100 -221 100
rect -163 -100 -93 100
rect -35 -100 35 100
rect 93 -100 163 100
rect 221 -100 291 100
rect 349 -100 419 100
rect 477 -100 547 100
<< pdiff >>
rect -605 88 -547 100
rect -605 -88 -593 88
rect -559 -88 -547 88
rect -605 -100 -547 -88
rect -477 88 -419 100
rect -477 -88 -465 88
rect -431 -88 -419 88
rect -477 -100 -419 -88
rect -349 88 -291 100
rect -349 -88 -337 88
rect -303 -88 -291 88
rect -349 -100 -291 -88
rect -221 88 -163 100
rect -221 -88 -209 88
rect -175 -88 -163 88
rect -221 -100 -163 -88
rect -93 88 -35 100
rect -93 -88 -81 88
rect -47 -88 -35 88
rect -93 -100 -35 -88
rect 35 88 93 100
rect 35 -88 47 88
rect 81 -88 93 88
rect 35 -100 93 -88
rect 163 88 221 100
rect 163 -88 175 88
rect 209 -88 221 88
rect 163 -100 221 -88
rect 291 88 349 100
rect 291 -88 303 88
rect 337 -88 349 88
rect 291 -100 349 -88
rect 419 88 477 100
rect 419 -88 431 88
rect 465 -88 477 88
rect 419 -100 477 -88
rect 547 88 605 100
rect 547 -88 559 88
rect 593 -88 605 88
rect 547 -100 605 -88
<< pdiffc >>
rect -593 -88 -559 88
rect -465 -88 -431 88
rect -337 -88 -303 88
rect -209 -88 -175 88
rect -81 -88 -47 88
rect 47 -88 81 88
rect 175 -88 209 88
rect 303 -88 337 88
rect 431 -88 465 88
rect 559 -88 593 88
<< nsubdiff >>
rect -707 276 -611 310
rect 611 276 707 310
rect -707 116 -673 276
rect 673 116 707 276
rect -707 -272 -673 -116
rect 673 -272 707 -116
rect -707 -306 -611 -272
rect 611 -306 707 -272
<< nsubdiffcont >>
rect -611 276 611 310
rect -707 -116 -673 116
rect 673 -116 707 116
rect -611 -306 611 -272
<< poly >>
rect -547 100 -477 126
rect -419 100 -349 126
rect -291 100 -221 126
rect -163 100 -93 126
rect -35 100 35 126
rect 93 100 163 126
rect 221 100 291 126
rect 349 100 419 126
rect 477 100 547 126
rect -547 -126 -477 -100
rect -419 -126 -349 -100
rect -291 -126 -221 -100
rect -163 -126 -93 -100
rect -35 -126 35 -100
rect 93 -126 163 -100
rect 221 -126 291 -100
rect 349 -126 419 -100
rect 477 -126 547 -100
<< locali >>
rect -707 276 -611 310
rect 611 276 707 310
rect -707 116 -673 276
rect 673 116 707 276
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -465 88 -431 104
rect -465 -104 -431 -88
rect -337 88 -303 104
rect -337 -104 -303 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -81 88 -47 104
rect -81 -104 -47 -88
rect 47 88 81 104
rect 47 -104 81 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 303 88 337 104
rect 303 -104 337 -88
rect 431 88 465 104
rect 431 -104 465 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect -707 -272 -673 -116
rect 673 -272 707 -116
rect -707 -306 -611 -272
rect 611 -306 707 -272
<< viali >>
rect -593 -88 -559 88
rect -465 -88 -431 88
rect -337 -88 -303 88
rect -209 -88 -175 88
rect -81 -88 -47 88
rect 47 -88 81 88
rect 175 -88 209 88
rect 303 -88 337 88
rect 431 -88 465 88
rect 559 -88 593 88
<< metal1 >>
rect -599 88 -553 100
rect -599 -88 -593 88
rect -559 -88 -553 88
rect -599 -100 -553 -88
rect -471 88 -425 100
rect -471 -88 -465 88
rect -431 -88 -425 88
rect -471 -100 -425 -88
rect -343 88 -297 100
rect -343 -88 -337 88
rect -303 -88 -297 88
rect -343 -100 -297 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -87 88 -41 100
rect -87 -88 -81 88
rect -47 -88 -41 88
rect -87 -100 -41 -88
rect 41 88 87 100
rect 41 -88 47 88
rect 81 -88 87 88
rect 41 -100 87 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 297 88 343 100
rect 297 -88 303 88
rect 337 -88 343 88
rect 297 -100 343 -88
rect 425 88 471 100
rect 425 -88 431 88
rect 465 -88 471 88
rect 425 -100 471 -88
rect 553 88 599 100
rect 553 -88 559 88
rect 593 -88 599 88
rect 553 -100 599 -88
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string FIXED_BBOX -690 -195 690 195
string parameters w 1 l 0.35 m 1 nf 9 diffcov 100 polycov 60 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1623971255
<< nwell >>
rect 9590 3318 13304 5174
rect 9590 -5978 13120 -4122
<< metal1 >>
rect 4664 -2760 4724 -2754
rect 4664 -3466 4724 -2820
rect 5690 -2822 5696 -2762
rect 5756 -2822 5762 -2762
rect 6602 -2822 6792 -2762
rect 5052 -3716 5112 -3398
rect 5308 -3716 5368 -3402
rect 5696 -3410 5756 -2822
rect 6080 -3716 6140 -3400
rect 6342 -3716 6402 -3404
rect 6732 -3414 6792 -2822
rect 16854 -3712 16914 -3430
rect 5046 -3776 5052 -3716
rect 5112 -3776 5118 -3716
rect 5302 -3776 5308 -3716
rect 5368 -3776 5374 -3716
rect 6074 -3776 6080 -3716
rect 6140 -3776 6146 -3716
rect 6336 -3776 6342 -3716
rect 6402 -3776 6408 -3716
rect 16848 -3772 16854 -3712
rect 16914 -3772 16920 -3712
<< via1 >>
rect 4664 -2820 4724 -2760
rect 5696 -2822 5756 -2762
rect 5052 -3776 5112 -3716
rect 5308 -3776 5368 -3716
rect 6080 -3776 6140 -3716
rect 6342 -3776 6402 -3716
rect 16854 -3772 16914 -3712
<< metal2 >>
rect 16973 3204 16982 3264
rect 17042 3204 17051 3264
rect 16982 3128 17042 3204
rect 4659 2928 4668 2988
rect 4728 2928 4737 2988
rect 11488 2871 11588 2876
rect 11484 2781 11493 2871
rect 11583 2781 11592 2871
rect 16459 2796 16468 2856
rect 16528 2796 17164 2856
rect 4998 2686 5184 2746
rect 9642 2740 9702 2749
rect 9578 2680 9642 2740
rect 9642 2671 9702 2680
rect 1489 1950 1498 2010
rect 1558 1950 1796 2010
rect 4732 1956 5170 2016
rect 6792 1050 6954 1110
rect 6772 -1914 6930 -1854
rect 4268 -2820 4664 -2760
rect 4724 -2820 4928 -2760
rect 5696 -2762 5756 -2756
rect 4268 -2916 4328 -2820
rect 5696 -2828 5756 -2822
rect 4259 -2976 4268 -2916
rect 4328 -2976 4337 -2916
rect 11488 -3464 11588 2781
rect 17734 2686 18144 2746
rect 18204 2686 18213 2746
rect 18156 1956 18980 2016
rect 11691 1816 11700 1916
rect 11800 1816 11809 1916
rect 11700 -2625 11800 1816
rect 18920 1684 18980 1956
rect 18911 1624 18920 1684
rect 18980 1624 18989 1684
rect 18536 1050 18740 1110
rect 18578 -1914 18742 -1854
rect 16979 -2462 16988 -2402
rect 17048 -2462 17057 -2402
rect 16988 -2522 17048 -2462
rect 16898 -2582 17048 -2522
rect 11696 -2715 11705 -2625
rect 11795 -2715 11804 -2625
rect 11700 -2720 11800 -2715
rect 16070 -2820 16720 -2760
rect 5045 -3550 5054 -3490
rect 5114 -3550 5304 -3490
rect 9286 -3544 9638 -3484
rect 9698 -3544 9707 -3484
rect 11479 -3564 11488 -3464
rect 11588 -3564 11597 -3464
rect 16070 -3480 16130 -2820
rect 16061 -3540 16070 -3480
rect 16130 -3540 16139 -3480
rect 21084 -3544 21440 -3484
rect 21500 -3544 21509 -3484
rect 5052 -3716 5112 -3710
rect 5308 -3716 5368 -3710
rect 6080 -3716 6140 -3710
rect 6342 -3716 6402 -3710
rect 16854 -3712 16914 -3706
rect 5112 -3776 5308 -3716
rect 5368 -3776 5492 -3716
rect 5980 -3776 6080 -3716
rect 6140 -3776 6342 -3716
rect 6402 -3776 6411 -3716
rect 16845 -3772 16854 -3712
rect 16914 -3772 16923 -3712
rect 5052 -3782 5112 -3776
rect 5308 -3782 5368 -3776
rect 6080 -3782 6140 -3776
rect 6342 -3782 6402 -3776
rect 16854 -3778 16914 -3772
<< via2 >>
rect 16982 3204 17042 3264
rect 4668 2928 4728 2988
rect 11493 2781 11583 2871
rect 16468 2796 16528 2856
rect 9642 2680 9702 2740
rect 1498 1950 1558 2010
rect 4268 -2976 4328 -2916
rect 18144 2686 18204 2746
rect 11700 1816 11800 1916
rect 18920 1624 18980 1684
rect 16988 -2462 17048 -2402
rect 11705 -2715 11795 -2625
rect 5054 -3550 5114 -3490
rect 9638 -3544 9698 -3484
rect 11488 -3564 11588 -3464
rect 16070 -3540 16130 -3480
rect 21440 -3544 21500 -3484
rect 6342 -3776 6402 -3716
rect 16854 -3772 16914 -3712
<< metal3 >>
rect 9620 3264 17070 3284
rect 9620 3204 16982 3264
rect 17042 3204 17070 3264
rect 9620 3184 17070 3204
rect -592 2988 4752 3008
rect -592 2928 4668 2988
rect 4728 2928 4752 2988
rect -592 2908 4752 2928
rect -592 -3466 -492 2908
rect 9620 2740 9720 3184
rect 11488 2871 16550 2876
rect 11488 2781 11493 2871
rect 11583 2856 16550 2871
rect 11583 2796 16468 2856
rect 16528 2796 16550 2856
rect 11583 2781 16550 2796
rect 11488 2776 16550 2781
rect 9620 2680 9642 2740
rect 9702 2680 9720 2740
rect 9620 2660 9720 2680
rect 18128 2746 23682 2764
rect 18128 2686 18144 2746
rect 18204 2686 23682 2746
rect 18128 2664 23682 2686
rect -330 2010 1580 2030
rect -330 1950 1498 2010
rect 1558 1950 1580 2010
rect -330 1930 1580 1950
rect -330 -2450 -230 1930
rect 11695 1916 11805 1921
rect 7896 1816 11700 1916
rect 11800 1816 16354 1916
rect 11695 1811 11805 1816
rect 18890 1684 23412 1706
rect 18890 1624 18920 1684
rect 18980 1624 23412 1684
rect 18890 1606 23412 1624
rect 23312 -2384 23412 1606
rect 16958 -2402 23412 -2384
rect -330 -2550 3908 -2450
rect 16958 -2462 16988 -2402
rect 17048 -2462 23412 -2402
rect 16958 -2484 23412 -2462
rect 3808 -2896 3908 -2550
rect 7972 -2625 16034 -2620
rect 7972 -2715 11705 -2625
rect 11795 -2715 16034 -2625
rect 7972 -2720 16034 -2715
rect 3808 -2916 4358 -2896
rect 3808 -2976 4268 -2916
rect 4328 -2976 4358 -2916
rect 3808 -2996 4358 -2976
rect 11483 -3464 11593 -3459
rect -592 -3490 5138 -3466
rect -592 -3550 5054 -3490
rect 5114 -3550 5138 -3490
rect -592 -3566 5138 -3550
rect 9614 -3484 11488 -3464
rect 9614 -3544 9638 -3484
rect 9698 -3544 11488 -3484
rect 9614 -3564 11488 -3544
rect 11588 -3480 16158 -3464
rect 23582 -3466 23682 2664
rect 11588 -3540 16070 -3480
rect 16130 -3540 16158 -3480
rect 11588 -3564 16158 -3540
rect 21422 -3484 23682 -3466
rect 21422 -3544 21440 -3484
rect 21500 -3544 23682 -3484
rect 11483 -3569 11593 -3564
rect 21422 -3566 23682 -3544
rect 6324 -3712 16934 -3696
rect 6324 -3716 16854 -3712
rect 6324 -3776 6342 -3716
rect 6402 -3772 16854 -3716
rect 16914 -3772 16934 -3712
rect 6402 -3776 16934 -3772
rect 6324 -3796 16934 -3776
<< metal4 >>
rect -728 4416 1572 5216
rect 9840 4416 12720 5216
rect 11292 -180 12036 434
rect -12 -624 23288 -180
rect 11292 -1242 12036 -624
rect -1528 -5246 1572 -5220
rect -1528 -5998 -1504 -5246
rect -752 -5998 1572 -5246
rect -1528 -6020 1572 -5998
rect 9904 -6020 12650 -5220
<< via4 >>
rect -1528 4416 -728 5216
rect -1504 -5998 -752 -5246
<< metal5 >>
rect -1552 5216 -704 5240
rect -1552 4416 -1528 5216
rect -728 4416 -704 5216
rect -1552 4392 -704 4416
rect -1528 -5246 -728 4392
rect -1528 -5998 -1504 -5246
rect -752 -5998 -728 -5246
rect -1528 -6022 -728 -5998
use gm_c_stage  gm_c_stage_2 gm_c_stage
timestamp 1623971255
transform 1 0 12188 0 1 2736
box -400 -3100 11100 2480
use gm_c_stage  gm_c_stage_3
timestamp 1623971255
transform 1 0 12188 0 -1 -3540
box -400 -3100 11100 2480
use gm_c_stage  gm_c_stage_1
timestamp 1623971255
transform 1 0 388 0 -1 -3540
box -400 -3100 11100 2480
use gm_c_stage  gm_c_stage_0
timestamp 1623971255
transform 1 0 388 0 1 2736
box -400 -3100 11100 2480
<< labels >>
flabel metal2 4746 1978 4762 1992 1 FreeSans 480 0 0 0 vip
flabel metal2 5012 2710 5020 2724 1 FreeSans 480 0 0 0 vim
flabel metal3 11604 1874 11614 1882 1 FreeSans 480 0 0 0 vocm
flabel metal4 11516 5188 11546 5206 1 FreeSans 480 0 0 0 VDD
flabel metal4 11416 -406 11440 -390 1 FreeSans 480 0 0 0 VSS
flabel metal3 23620 1100 23640 1116 1 FreeSans 480 0 0 0 vfiltm
flabel metal3 23360 1060 23382 1076 1 FreeSans 480 0 0 0 vfiltp
flabel metal3 -562 1138 -542 1158 1 FreeSans 480 0 0 0 vintp
flabel metal3 -290 1124 -268 1144 1 FreeSans 480 0 0 0 vintm
flabel metal2 6858 1072 6874 1080 1 FreeSans 480 0 0 0 ibiasn1
flabel metal2 6844 -1890 6870 -1878 1 FreeSans 480 0 0 0 ibiasn2
flabel metal2 18656 -1896 18670 -1880 1 FreeSans 480 0 0 0 ibiasn3
flabel metal2 18640 1074 18656 1084 1 FreeSans 480 0 0 0 ibiasn4
<< end >>
